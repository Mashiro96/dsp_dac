module DspDecode(
  input         clock,
  input         reset,
  output        io_din_ready,
  input         io_din_valid,
  input  [31:0] io_din_bits_0,
  input  [31:0] io_din_bits_1,
  input         io_dout_ready,
  output        io_dout_valid,
  output [31:0] io_dout_bits_0,
  output [31:0] io_dout_bits_1,
  input         io_macuio_0_ready,
  output        io_macuio_0_valid,
  output [2:0]  io_macuio_0_bits_vlen,
  output        io_macuio_0_bits_select,
  output        io_macuio_0_bits_drc,
  output        io_macuio_0_bits_pow,
  output        io_macuio_0_bits_loop,
  output        io_macuio_0_bits_drcgain,
  output        io_macuio_0_bits_drcnum,
  output        io_macuio_0_bits_srcreq_0_valid,
  output        io_macuio_0_bits_srcreq_0_isgroup,
  output        io_macuio_0_bits_srcreq_0_iscoef,
  output [5:0]  io_macuio_0_bits_srcreq_0_idx,
  output        io_macuio_0_bits_srcreq_0_busy,
  output        io_macuio_0_bits_srcreq_0_wkupidx_0,
  output        io_macuio_0_bits_srcreq_0_wkupidx_1,
  output        io_macuio_0_bits_srcreq_0_wkupidx_2,
  output        io_macuio_0_bits_srcreq_0_wkupidx_3,
  output        io_macuio_0_bits_srcreq_0_wkupidx_4,
  output        io_macuio_0_bits_srcreq_0_wkupidx_5,
  output        io_macuio_0_bits_srcreq_1_valid,
  output        io_macuio_0_bits_srcreq_1_isgroup,
  output        io_macuio_0_bits_srcreq_1_iscoef,
  output [5:0]  io_macuio_0_bits_srcreq_1_idx,
  output        io_macuio_0_bits_srcreq_1_busy,
  output        io_macuio_0_bits_srcreq_1_wkupidx_0,
  output        io_macuio_0_bits_srcreq_1_wkupidx_1,
  output        io_macuio_0_bits_srcreq_1_wkupidx_2,
  output        io_macuio_0_bits_srcreq_1_wkupidx_3,
  output        io_macuio_0_bits_srcreq_1_wkupidx_4,
  output        io_macuio_0_bits_srcreq_1_wkupidx_5,
  output        io_macuio_0_bits_srcreq_2_valid,
  output        io_macuio_0_bits_srcreq_2_isgroup,
  output        io_macuio_0_bits_srcreq_2_iscoef,
  output [5:0]  io_macuio_0_bits_srcreq_2_idx,
  output        io_macuio_0_bits_srcreq_2_busy,
  output        io_macuio_0_bits_srcreq_2_wkupidx_0,
  output        io_macuio_0_bits_srcreq_2_wkupidx_1,
  output        io_macuio_0_bits_srcreq_2_wkupidx_2,
  output        io_macuio_0_bits_srcreq_2_wkupidx_3,
  output        io_macuio_0_bits_srcreq_2_wkupidx_4,
  output        io_macuio_0_bits_srcreq_2_wkupidx_5,
  output        io_macuio_0_bits_srcreq_3_valid,
  output        io_macuio_0_bits_srcreq_3_isgroup,
  output        io_macuio_0_bits_srcreq_3_iscoef,
  output [5:0]  io_macuio_0_bits_srcreq_3_idx,
  output        io_macuio_0_bits_srcreq_3_busy,
  output        io_macuio_0_bits_srcreq_3_wkupidx_0,
  output        io_macuio_0_bits_srcreq_3_wkupidx_1,
  output        io_macuio_0_bits_srcreq_3_wkupidx_2,
  output        io_macuio_0_bits_srcreq_3_wkupidx_3,
  output        io_macuio_0_bits_srcreq_3_wkupidx_4,
  output        io_macuio_0_bits_srcreq_3_wkupidx_5,
  output        io_macuio_0_bits_srcreq_4_valid,
  output        io_macuio_0_bits_srcreq_4_isgroup,
  output        io_macuio_0_bits_srcreq_4_iscoef,
  output [5:0]  io_macuio_0_bits_srcreq_4_idx,
  output        io_macuio_0_bits_srcreq_4_busy,
  output        io_macuio_0_bits_srcreq_4_wkupidx_0,
  output        io_macuio_0_bits_srcreq_4_wkupidx_1,
  output        io_macuio_0_bits_srcreq_4_wkupidx_2,
  output        io_macuio_0_bits_srcreq_4_wkupidx_3,
  output        io_macuio_0_bits_srcreq_4_wkupidx_4,
  output        io_macuio_0_bits_srcreq_4_wkupidx_5,
  output        io_macuio_0_bits_srcreq_5_valid,
  output        io_macuio_0_bits_srcreq_5_isgroup,
  output        io_macuio_0_bits_srcreq_5_iscoef,
  output [5:0]  io_macuio_0_bits_srcreq_5_idx,
  output        io_macuio_0_bits_srcreq_5_busy,
  output        io_macuio_0_bits_srcreq_5_wkupidx_0,
  output        io_macuio_0_bits_srcreq_5_wkupidx_1,
  output        io_macuio_0_bits_srcreq_5_wkupidx_2,
  output        io_macuio_0_bits_srcreq_5_wkupidx_3,
  output        io_macuio_0_bits_srcreq_5_wkupidx_4,
  output        io_macuio_0_bits_srcreq_5_wkupidx_5,
  output        io_macuio_0_bits_wbvld,
  output [5:0]  io_macuio_0_bits_wbreq,
  output        io_macuio_0_bits_waridx_0,
  output        io_macuio_0_bits_waridx_1,
  output        io_macuio_0_bits_waridx_2,
  output        io_macuio_0_bits_waridx_3,
  output        io_macuio_0_bits_waridx_4,
  output        io_macuio_0_bits_wawidx_0,
  output        io_macuio_0_bits_wawidx_1,
  output        io_macuio_0_bits_wawidx_2,
  output        io_macuio_0_bits_wawidx_3,
  output        io_macuio_0_bits_wawidx_4,
  input         io_macuio_1_ready,
  output        io_macuio_1_valid,
  output [2:0]  io_macuio_1_bits_vlen,
  output        io_macuio_1_bits_select,
  output        io_macuio_1_bits_drc,
  output        io_macuio_1_bits_pow,
  output        io_macuio_1_bits_loop,
  output        io_macuio_1_bits_drcgain,
  output        io_macuio_1_bits_drcnum,
  output        io_macuio_1_bits_srcreq_0_valid,
  output        io_macuio_1_bits_srcreq_0_isgroup,
  output        io_macuio_1_bits_srcreq_0_iscoef,
  output [5:0]  io_macuio_1_bits_srcreq_0_idx,
  output        io_macuio_1_bits_srcreq_0_busy,
  output        io_macuio_1_bits_srcreq_0_wkupidx_0,
  output        io_macuio_1_bits_srcreq_0_wkupidx_1,
  output        io_macuio_1_bits_srcreq_0_wkupidx_2,
  output        io_macuio_1_bits_srcreq_0_wkupidx_3,
  output        io_macuio_1_bits_srcreq_0_wkupidx_4,
  output        io_macuio_1_bits_srcreq_0_wkupidx_5,
  output        io_macuio_1_bits_srcreq_1_valid,
  output        io_macuio_1_bits_srcreq_1_isgroup,
  output        io_macuio_1_bits_srcreq_1_iscoef,
  output [5:0]  io_macuio_1_bits_srcreq_1_idx,
  output        io_macuio_1_bits_srcreq_1_busy,
  output        io_macuio_1_bits_srcreq_1_wkupidx_0,
  output        io_macuio_1_bits_srcreq_1_wkupidx_1,
  output        io_macuio_1_bits_srcreq_1_wkupidx_2,
  output        io_macuio_1_bits_srcreq_1_wkupidx_3,
  output        io_macuio_1_bits_srcreq_1_wkupidx_4,
  output        io_macuio_1_bits_srcreq_1_wkupidx_5,
  output        io_macuio_1_bits_srcreq_2_valid,
  output        io_macuio_1_bits_srcreq_2_isgroup,
  output        io_macuio_1_bits_srcreq_2_iscoef,
  output [5:0]  io_macuio_1_bits_srcreq_2_idx,
  output        io_macuio_1_bits_srcreq_2_busy,
  output        io_macuio_1_bits_srcreq_2_wkupidx_0,
  output        io_macuio_1_bits_srcreq_2_wkupidx_1,
  output        io_macuio_1_bits_srcreq_2_wkupidx_2,
  output        io_macuio_1_bits_srcreq_2_wkupidx_3,
  output        io_macuio_1_bits_srcreq_2_wkupidx_4,
  output        io_macuio_1_bits_srcreq_2_wkupidx_5,
  output        io_macuio_1_bits_srcreq_3_valid,
  output        io_macuio_1_bits_srcreq_3_isgroup,
  output        io_macuio_1_bits_srcreq_3_iscoef,
  output [5:0]  io_macuio_1_bits_srcreq_3_idx,
  output        io_macuio_1_bits_srcreq_3_busy,
  output        io_macuio_1_bits_srcreq_3_wkupidx_0,
  output        io_macuio_1_bits_srcreq_3_wkupidx_1,
  output        io_macuio_1_bits_srcreq_3_wkupidx_2,
  output        io_macuio_1_bits_srcreq_3_wkupidx_3,
  output        io_macuio_1_bits_srcreq_3_wkupidx_4,
  output        io_macuio_1_bits_srcreq_3_wkupidx_5,
  output        io_macuio_1_bits_srcreq_4_valid,
  output        io_macuio_1_bits_srcreq_4_isgroup,
  output        io_macuio_1_bits_srcreq_4_iscoef,
  output [5:0]  io_macuio_1_bits_srcreq_4_idx,
  output        io_macuio_1_bits_srcreq_4_busy,
  output        io_macuio_1_bits_srcreq_4_wkupidx_0,
  output        io_macuio_1_bits_srcreq_4_wkupidx_1,
  output        io_macuio_1_bits_srcreq_4_wkupidx_2,
  output        io_macuio_1_bits_srcreq_4_wkupidx_3,
  output        io_macuio_1_bits_srcreq_4_wkupidx_4,
  output        io_macuio_1_bits_srcreq_4_wkupidx_5,
  output        io_macuio_1_bits_srcreq_5_valid,
  output        io_macuio_1_bits_srcreq_5_isgroup,
  output        io_macuio_1_bits_srcreq_5_iscoef,
  output [5:0]  io_macuio_1_bits_srcreq_5_idx,
  output        io_macuio_1_bits_srcreq_5_busy,
  output        io_macuio_1_bits_srcreq_5_wkupidx_0,
  output        io_macuio_1_bits_srcreq_5_wkupidx_1,
  output        io_macuio_1_bits_srcreq_5_wkupidx_2,
  output        io_macuio_1_bits_srcreq_5_wkupidx_3,
  output        io_macuio_1_bits_srcreq_5_wkupidx_4,
  output        io_macuio_1_bits_srcreq_5_wkupidx_5,
  output        io_macuio_1_bits_wbvld,
  output [5:0]  io_macuio_1_bits_wbreq,
  output        io_macuio_1_bits_waridx_0,
  output        io_macuio_1_bits_waridx_1,
  output        io_macuio_1_bits_waridx_2,
  output        io_macuio_1_bits_waridx_3,
  output        io_macuio_1_bits_waridx_4,
  output        io_macuio_1_bits_wawidx_0,
  output        io_macuio_1_bits_wawidx_1,
  output        io_macuio_1_bits_wawidx_2,
  output        io_macuio_1_bits_wawidx_3,
  output        io_macuio_1_bits_wawidx_4,
  input         io_macuio_2_ready,
  output        io_macuio_2_valid,
  output [2:0]  io_macuio_2_bits_vlen,
  output        io_macuio_2_bits_select,
  output        io_macuio_2_bits_drc,
  output        io_macuio_2_bits_pow,
  output        io_macuio_2_bits_loop,
  output        io_macuio_2_bits_drcgain,
  output        io_macuio_2_bits_drcnum,
  output        io_macuio_2_bits_srcreq_0_valid,
  output        io_macuio_2_bits_srcreq_0_isgroup,
  output        io_macuio_2_bits_srcreq_0_iscoef,
  output [5:0]  io_macuio_2_bits_srcreq_0_idx,
  output        io_macuio_2_bits_srcreq_0_busy,
  output        io_macuio_2_bits_srcreq_0_wkupidx_0,
  output        io_macuio_2_bits_srcreq_0_wkupidx_1,
  output        io_macuio_2_bits_srcreq_0_wkupidx_2,
  output        io_macuio_2_bits_srcreq_0_wkupidx_3,
  output        io_macuio_2_bits_srcreq_0_wkupidx_4,
  output        io_macuio_2_bits_srcreq_0_wkupidx_5,
  output        io_macuio_2_bits_srcreq_1_valid,
  output        io_macuio_2_bits_srcreq_1_isgroup,
  output        io_macuio_2_bits_srcreq_1_iscoef,
  output [5:0]  io_macuio_2_bits_srcreq_1_idx,
  output        io_macuio_2_bits_srcreq_1_busy,
  output        io_macuio_2_bits_srcreq_1_wkupidx_0,
  output        io_macuio_2_bits_srcreq_1_wkupidx_1,
  output        io_macuio_2_bits_srcreq_1_wkupidx_2,
  output        io_macuio_2_bits_srcreq_1_wkupidx_3,
  output        io_macuio_2_bits_srcreq_1_wkupidx_4,
  output        io_macuio_2_bits_srcreq_1_wkupidx_5,
  output        io_macuio_2_bits_srcreq_2_valid,
  output        io_macuio_2_bits_srcreq_2_isgroup,
  output        io_macuio_2_bits_srcreq_2_iscoef,
  output [5:0]  io_macuio_2_bits_srcreq_2_idx,
  output        io_macuio_2_bits_srcreq_2_busy,
  output        io_macuio_2_bits_srcreq_2_wkupidx_0,
  output        io_macuio_2_bits_srcreq_2_wkupidx_1,
  output        io_macuio_2_bits_srcreq_2_wkupidx_2,
  output        io_macuio_2_bits_srcreq_2_wkupidx_3,
  output        io_macuio_2_bits_srcreq_2_wkupidx_4,
  output        io_macuio_2_bits_srcreq_2_wkupidx_5,
  output        io_macuio_2_bits_srcreq_3_valid,
  output        io_macuio_2_bits_srcreq_3_isgroup,
  output        io_macuio_2_bits_srcreq_3_iscoef,
  output [5:0]  io_macuio_2_bits_srcreq_3_idx,
  output        io_macuio_2_bits_srcreq_3_busy,
  output        io_macuio_2_bits_srcreq_3_wkupidx_0,
  output        io_macuio_2_bits_srcreq_3_wkupidx_1,
  output        io_macuio_2_bits_srcreq_3_wkupidx_2,
  output        io_macuio_2_bits_srcreq_3_wkupidx_3,
  output        io_macuio_2_bits_srcreq_3_wkupidx_4,
  output        io_macuio_2_bits_srcreq_3_wkupidx_5,
  output        io_macuio_2_bits_srcreq_4_valid,
  output        io_macuio_2_bits_srcreq_4_isgroup,
  output        io_macuio_2_bits_srcreq_4_iscoef,
  output [5:0]  io_macuio_2_bits_srcreq_4_idx,
  output        io_macuio_2_bits_srcreq_4_busy,
  output        io_macuio_2_bits_srcreq_4_wkupidx_0,
  output        io_macuio_2_bits_srcreq_4_wkupidx_1,
  output        io_macuio_2_bits_srcreq_4_wkupidx_2,
  output        io_macuio_2_bits_srcreq_4_wkupidx_3,
  output        io_macuio_2_bits_srcreq_4_wkupidx_4,
  output        io_macuio_2_bits_srcreq_4_wkupidx_5,
  output        io_macuio_2_bits_srcreq_5_valid,
  output        io_macuio_2_bits_srcreq_5_isgroup,
  output        io_macuio_2_bits_srcreq_5_iscoef,
  output [5:0]  io_macuio_2_bits_srcreq_5_idx,
  output        io_macuio_2_bits_srcreq_5_busy,
  output        io_macuio_2_bits_srcreq_5_wkupidx_0,
  output        io_macuio_2_bits_srcreq_5_wkupidx_1,
  output        io_macuio_2_bits_srcreq_5_wkupidx_2,
  output        io_macuio_2_bits_srcreq_5_wkupidx_3,
  output        io_macuio_2_bits_srcreq_5_wkupidx_4,
  output        io_macuio_2_bits_srcreq_5_wkupidx_5,
  output        io_macuio_2_bits_wbvld,
  output [5:0]  io_macuio_2_bits_wbreq,
  output        io_macuio_2_bits_waridx_0,
  output        io_macuio_2_bits_waridx_1,
  output        io_macuio_2_bits_waridx_2,
  output        io_macuio_2_bits_waridx_3,
  output        io_macuio_2_bits_waridx_4,
  output        io_macuio_2_bits_wawidx_0,
  output        io_macuio_2_bits_wawidx_1,
  output        io_macuio_2_bits_wawidx_2,
  output        io_macuio_2_bits_wawidx_3,
  output        io_macuio_2_bits_wawidx_4,
  input         io_macuio_3_ready,
  output        io_macuio_3_valid,
  output [2:0]  io_macuio_3_bits_vlen,
  output        io_macuio_3_bits_select,
  output        io_macuio_3_bits_drc,
  output        io_macuio_3_bits_pow,
  output        io_macuio_3_bits_loop,
  output        io_macuio_3_bits_drcgain,
  output        io_macuio_3_bits_drcnum,
  output        io_macuio_3_bits_srcreq_0_valid,
  output        io_macuio_3_bits_srcreq_0_isgroup,
  output        io_macuio_3_bits_srcreq_0_iscoef,
  output [5:0]  io_macuio_3_bits_srcreq_0_idx,
  output        io_macuio_3_bits_srcreq_0_busy,
  output        io_macuio_3_bits_srcreq_0_wkupidx_0,
  output        io_macuio_3_bits_srcreq_0_wkupidx_1,
  output        io_macuio_3_bits_srcreq_0_wkupidx_2,
  output        io_macuio_3_bits_srcreq_0_wkupidx_3,
  output        io_macuio_3_bits_srcreq_0_wkupidx_4,
  output        io_macuio_3_bits_srcreq_0_wkupidx_5,
  output        io_macuio_3_bits_srcreq_1_valid,
  output        io_macuio_3_bits_srcreq_1_isgroup,
  output        io_macuio_3_bits_srcreq_1_iscoef,
  output [5:0]  io_macuio_3_bits_srcreq_1_idx,
  output        io_macuio_3_bits_srcreq_1_busy,
  output        io_macuio_3_bits_srcreq_1_wkupidx_0,
  output        io_macuio_3_bits_srcreq_1_wkupidx_1,
  output        io_macuio_3_bits_srcreq_1_wkupidx_2,
  output        io_macuio_3_bits_srcreq_1_wkupidx_3,
  output        io_macuio_3_bits_srcreq_1_wkupidx_4,
  output        io_macuio_3_bits_srcreq_1_wkupidx_5,
  output        io_macuio_3_bits_srcreq_2_valid,
  output        io_macuio_3_bits_srcreq_2_isgroup,
  output        io_macuio_3_bits_srcreq_2_iscoef,
  output [5:0]  io_macuio_3_bits_srcreq_2_idx,
  output        io_macuio_3_bits_srcreq_2_busy,
  output        io_macuio_3_bits_srcreq_2_wkupidx_0,
  output        io_macuio_3_bits_srcreq_2_wkupidx_1,
  output        io_macuio_3_bits_srcreq_2_wkupidx_2,
  output        io_macuio_3_bits_srcreq_2_wkupidx_3,
  output        io_macuio_3_bits_srcreq_2_wkupidx_4,
  output        io_macuio_3_bits_srcreq_2_wkupidx_5,
  output        io_macuio_3_bits_srcreq_3_valid,
  output        io_macuio_3_bits_srcreq_3_isgroup,
  output        io_macuio_3_bits_srcreq_3_iscoef,
  output [5:0]  io_macuio_3_bits_srcreq_3_idx,
  output        io_macuio_3_bits_srcreq_3_busy,
  output        io_macuio_3_bits_srcreq_3_wkupidx_0,
  output        io_macuio_3_bits_srcreq_3_wkupidx_1,
  output        io_macuio_3_bits_srcreq_3_wkupidx_2,
  output        io_macuio_3_bits_srcreq_3_wkupidx_3,
  output        io_macuio_3_bits_srcreq_3_wkupidx_4,
  output        io_macuio_3_bits_srcreq_3_wkupidx_5,
  output        io_macuio_3_bits_srcreq_4_valid,
  output        io_macuio_3_bits_srcreq_4_isgroup,
  output        io_macuio_3_bits_srcreq_4_iscoef,
  output [5:0]  io_macuio_3_bits_srcreq_4_idx,
  output        io_macuio_3_bits_srcreq_4_busy,
  output        io_macuio_3_bits_srcreq_4_wkupidx_0,
  output        io_macuio_3_bits_srcreq_4_wkupidx_1,
  output        io_macuio_3_bits_srcreq_4_wkupidx_2,
  output        io_macuio_3_bits_srcreq_4_wkupidx_3,
  output        io_macuio_3_bits_srcreq_4_wkupidx_4,
  output        io_macuio_3_bits_srcreq_4_wkupidx_5,
  output        io_macuio_3_bits_srcreq_5_valid,
  output        io_macuio_3_bits_srcreq_5_isgroup,
  output        io_macuio_3_bits_srcreq_5_iscoef,
  output [5:0]  io_macuio_3_bits_srcreq_5_idx,
  output        io_macuio_3_bits_srcreq_5_busy,
  output        io_macuio_3_bits_srcreq_5_wkupidx_0,
  output        io_macuio_3_bits_srcreq_5_wkupidx_1,
  output        io_macuio_3_bits_srcreq_5_wkupidx_2,
  output        io_macuio_3_bits_srcreq_5_wkupidx_3,
  output        io_macuio_3_bits_srcreq_5_wkupidx_4,
  output        io_macuio_3_bits_srcreq_5_wkupidx_5,
  output        io_macuio_3_bits_wbvld,
  output [5:0]  io_macuio_3_bits_wbreq,
  output        io_macuio_3_bits_waridx_0,
  output        io_macuio_3_bits_waridx_1,
  output        io_macuio_3_bits_waridx_2,
  output        io_macuio_3_bits_waridx_3,
  output        io_macuio_3_bits_waridx_4,
  output        io_macuio_3_bits_wawidx_0,
  output        io_macuio_3_bits_wawidx_1,
  output        io_macuio_3_bits_wawidx_2,
  output        io_macuio_3_bits_wawidx_3,
  output        io_macuio_3_bits_wawidx_4,
  input         io_macuio_4_ready,
  output        io_macuio_4_valid,
  output [2:0]  io_macuio_4_bits_vlen,
  output        io_macuio_4_bits_select,
  output        io_macuio_4_bits_drc,
  output        io_macuio_4_bits_pow,
  output        io_macuio_4_bits_loop,
  output        io_macuio_4_bits_drcgain,
  output        io_macuio_4_bits_drcnum,
  output        io_macuio_4_bits_srcreq_0_valid,
  output        io_macuio_4_bits_srcreq_0_isgroup,
  output        io_macuio_4_bits_srcreq_0_iscoef,
  output [5:0]  io_macuio_4_bits_srcreq_0_idx,
  output        io_macuio_4_bits_srcreq_0_busy,
  output        io_macuio_4_bits_srcreq_0_wkupidx_0,
  output        io_macuio_4_bits_srcreq_0_wkupidx_1,
  output        io_macuio_4_bits_srcreq_0_wkupidx_2,
  output        io_macuio_4_bits_srcreq_0_wkupidx_3,
  output        io_macuio_4_bits_srcreq_0_wkupidx_4,
  output        io_macuio_4_bits_srcreq_0_wkupidx_5,
  output        io_macuio_4_bits_srcreq_1_valid,
  output        io_macuio_4_bits_srcreq_1_isgroup,
  output        io_macuio_4_bits_srcreq_1_iscoef,
  output [5:0]  io_macuio_4_bits_srcreq_1_idx,
  output        io_macuio_4_bits_srcreq_1_busy,
  output        io_macuio_4_bits_srcreq_1_wkupidx_0,
  output        io_macuio_4_bits_srcreq_1_wkupidx_1,
  output        io_macuio_4_bits_srcreq_1_wkupidx_2,
  output        io_macuio_4_bits_srcreq_1_wkupidx_3,
  output        io_macuio_4_bits_srcreq_1_wkupidx_4,
  output        io_macuio_4_bits_srcreq_1_wkupidx_5,
  output        io_macuio_4_bits_srcreq_2_valid,
  output        io_macuio_4_bits_srcreq_2_isgroup,
  output        io_macuio_4_bits_srcreq_2_iscoef,
  output [5:0]  io_macuio_4_bits_srcreq_2_idx,
  output        io_macuio_4_bits_srcreq_2_busy,
  output        io_macuio_4_bits_srcreq_2_wkupidx_0,
  output        io_macuio_4_bits_srcreq_2_wkupidx_1,
  output        io_macuio_4_bits_srcreq_2_wkupidx_2,
  output        io_macuio_4_bits_srcreq_2_wkupidx_3,
  output        io_macuio_4_bits_srcreq_2_wkupidx_4,
  output        io_macuio_4_bits_srcreq_2_wkupidx_5,
  output        io_macuio_4_bits_srcreq_3_valid,
  output        io_macuio_4_bits_srcreq_3_isgroup,
  output        io_macuio_4_bits_srcreq_3_iscoef,
  output [5:0]  io_macuio_4_bits_srcreq_3_idx,
  output        io_macuio_4_bits_srcreq_3_busy,
  output        io_macuio_4_bits_srcreq_3_wkupidx_0,
  output        io_macuio_4_bits_srcreq_3_wkupidx_1,
  output        io_macuio_4_bits_srcreq_3_wkupidx_2,
  output        io_macuio_4_bits_srcreq_3_wkupidx_3,
  output        io_macuio_4_bits_srcreq_3_wkupidx_4,
  output        io_macuio_4_bits_srcreq_3_wkupidx_5,
  output        io_macuio_4_bits_srcreq_4_valid,
  output        io_macuio_4_bits_srcreq_4_isgroup,
  output        io_macuio_4_bits_srcreq_4_iscoef,
  output [5:0]  io_macuio_4_bits_srcreq_4_idx,
  output        io_macuio_4_bits_srcreq_4_busy,
  output        io_macuio_4_bits_srcreq_4_wkupidx_0,
  output        io_macuio_4_bits_srcreq_4_wkupidx_1,
  output        io_macuio_4_bits_srcreq_4_wkupidx_2,
  output        io_macuio_4_bits_srcreq_4_wkupidx_3,
  output        io_macuio_4_bits_srcreq_4_wkupidx_4,
  output        io_macuio_4_bits_srcreq_4_wkupidx_5,
  output        io_macuio_4_bits_srcreq_5_valid,
  output        io_macuio_4_bits_srcreq_5_isgroup,
  output        io_macuio_4_bits_srcreq_5_iscoef,
  output [5:0]  io_macuio_4_bits_srcreq_5_idx,
  output        io_macuio_4_bits_srcreq_5_busy,
  output        io_macuio_4_bits_srcreq_5_wkupidx_0,
  output        io_macuio_4_bits_srcreq_5_wkupidx_1,
  output        io_macuio_4_bits_srcreq_5_wkupidx_2,
  output        io_macuio_4_bits_srcreq_5_wkupidx_3,
  output        io_macuio_4_bits_srcreq_5_wkupidx_4,
  output        io_macuio_4_bits_srcreq_5_wkupidx_5,
  output        io_macuio_4_bits_wbvld,
  output [5:0]  io_macuio_4_bits_wbreq,
  output        io_macuio_4_bits_waridx_0,
  output        io_macuio_4_bits_waridx_1,
  output        io_macuio_4_bits_waridx_2,
  output        io_macuio_4_bits_waridx_3,
  output        io_macuio_4_bits_waridx_4,
  output        io_macuio_4_bits_wawidx_0,
  output        io_macuio_4_bits_wawidx_1,
  output        io_macuio_4_bits_wawidx_2,
  output        io_macuio_4_bits_wawidx_3,
  output        io_macuio_4_bits_wawidx_4,
  input         io_wd_check_0_valid,
  input  [5:0]  io_wd_check_0_bits,
  input         io_wd_check_1_valid,
  input  [5:0]  io_wd_check_1_bits,
  input         io_wd_check_2_valid,
  input  [5:0]  io_wd_check_2_bits,
  input         io_wd_check_3_valid,
  input  [5:0]  io_wd_check_3_bits,
  input         io_wd_check_4_valid,
  input  [5:0]  io_wd_check_4_bits,
  input         io_wd_check_5_valid,
  input  [5:0]  io_wd_check_5_bits,
  input         io_mac_r_check_0_0_valid,
  input  [5:0]  io_mac_r_check_0_0_bits,
  input         io_mac_r_check_0_1_valid,
  input  [5:0]  io_mac_r_check_0_1_bits,
  input         io_mac_r_check_0_2_valid,
  input  [5:0]  io_mac_r_check_0_2_bits,
  input         io_mac_r_check_0_3_valid,
  input  [5:0]  io_mac_r_check_0_3_bits,
  input         io_mac_r_check_0_4_valid,
  input  [5:0]  io_mac_r_check_0_4_bits,
  input         io_mac_r_check_0_5_valid,
  input  [5:0]  io_mac_r_check_0_5_bits,
  input         io_mac_r_check_1_0_valid,
  input  [5:0]  io_mac_r_check_1_0_bits,
  input         io_mac_r_check_1_1_valid,
  input  [5:0]  io_mac_r_check_1_1_bits,
  input         io_mac_r_check_1_2_valid,
  input  [5:0]  io_mac_r_check_1_2_bits,
  input         io_mac_r_check_1_3_valid,
  input  [5:0]  io_mac_r_check_1_3_bits,
  input         io_mac_r_check_1_4_valid,
  input  [5:0]  io_mac_r_check_1_4_bits,
  input         io_mac_r_check_1_5_valid,
  input  [5:0]  io_mac_r_check_1_5_bits,
  input         io_mac_r_check_2_0_valid,
  input  [5:0]  io_mac_r_check_2_0_bits,
  input         io_mac_r_check_2_1_valid,
  input  [5:0]  io_mac_r_check_2_1_bits,
  input         io_mac_r_check_2_2_valid,
  input  [5:0]  io_mac_r_check_2_2_bits,
  input         io_mac_r_check_2_3_valid,
  input  [5:0]  io_mac_r_check_2_3_bits,
  input         io_mac_r_check_2_4_valid,
  input  [5:0]  io_mac_r_check_2_4_bits,
  input         io_mac_r_check_2_5_valid,
  input  [5:0]  io_mac_r_check_2_5_bits,
  input         io_mac_r_check_3_0_valid,
  input  [5:0]  io_mac_r_check_3_0_bits,
  input         io_mac_r_check_3_1_valid,
  input  [5:0]  io_mac_r_check_3_1_bits,
  input         io_mac_r_check_3_2_valid,
  input  [5:0]  io_mac_r_check_3_2_bits,
  input         io_mac_r_check_3_3_valid,
  input  [5:0]  io_mac_r_check_3_3_bits,
  input         io_mac_r_check_3_4_valid,
  input  [5:0]  io_mac_r_check_3_4_bits,
  input         io_mac_r_check_3_5_valid,
  input  [5:0]  io_mac_r_check_3_5_bits,
  input         io_mac_r_check_4_0_valid,
  input  [5:0]  io_mac_r_check_4_0_bits,
  input         io_mac_r_check_4_1_valid,
  input  [5:0]  io_mac_r_check_4_1_bits,
  input         io_mac_r_check_4_2_valid,
  input  [5:0]  io_mac_r_check_4_2_bits,
  input         io_mac_r_check_4_3_valid,
  input  [5:0]  io_mac_r_check_4_3_bits,
  input         io_mac_r_check_4_4_valid,
  input  [5:0]  io_mac_r_check_4_4_bits,
  input         io_mac_r_check_4_5_valid,
  input  [5:0]  io_mac_r_check_4_5_bits,
  input         io_cor_r_check_0_valid,
  input  [5:0]  io_cor_r_check_0_bits,
  input         io_cor_r_check_1_valid,
  input  [5:0]  io_cor_r_check_1_bits,
  input         io_exuempty_0,
  input         io_exuempty_1,
  input         io_exuempty_2,
  input         io_exuempty_3,
  input         io_exuempty_4,
  input         io_exuempty_5,
  input         io_coruio_ready,
  output        io_coruio_valid,
  output        io_coruio_bits_cortype,
  output        io_coruio_bits_srcreq_0_valid,
  output [5:0]  io_coruio_bits_srcreq_0_idx,
  output        io_coruio_bits_srcreq_0_busy,
  output        io_coruio_bits_srcreq_0_wkupidx_0,
  output        io_coruio_bits_srcreq_0_wkupidx_1,
  output        io_coruio_bits_srcreq_0_wkupidx_2,
  output        io_coruio_bits_srcreq_0_wkupidx_3,
  output        io_coruio_bits_srcreq_0_wkupidx_4,
  output        io_coruio_bits_srcreq_0_wkupidx_5,
  output        io_coruio_bits_srcreq_1_valid,
  output [5:0]  io_coruio_bits_srcreq_1_idx,
  output        io_coruio_bits_srcreq_1_busy,
  output        io_coruio_bits_srcreq_1_wkupidx_0,
  output        io_coruio_bits_srcreq_1_wkupidx_1,
  output        io_coruio_bits_srcreq_1_wkupidx_2,
  output        io_coruio_bits_srcreq_1_wkupidx_3,
  output        io_coruio_bits_srcreq_1_wkupidx_4,
  output        io_coruio_bits_srcreq_1_wkupidx_5,
  output        io_coruio_bits_wbvld,
  output [5:0]  io_coruio_bits_wbreq,
  output        io_coruio_bits_waridx_0,
  output        io_coruio_bits_waridx_1,
  output        io_coruio_bits_waridx_2,
  output        io_coruio_bits_waridx_3,
  output        io_coruio_bits_waridx_4,
  output        io_coruio_bits_wawidx_0,
  output        io_coruio_bits_wawidx_1,
  output        io_coruio_bits_wawidx_2,
  output        io_coruio_bits_wawidx_3,
  output        io_coruio_bits_wawidx_4,
  output        io_writerf_valid,
  output [31:0] io_writerf_bits_0,
  output [31:0] io_writerf_bits_1,
  output [31:0] io_writerf_bits_2,
  output [31:0] io_writerf_bits_3,
  input  [31:0] io_readrf_0,
  input  [31:0] io_readrf_1,
  input  [2:0]  io_coef_in_mainch_ch0_inputsel,
  input  [2:0]  io_coef_in_mainch_ch1_inputsel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] instcnt; // @[dspdecode.scala 75:24]
  wire [8:0] _GEN_1 = 6'h1 == instcnt ? 9'h2 : 9'h0; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_2 = 6'h2 == instcnt ? 9'h52 : _GEN_1; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_3 = 6'h3 == instcnt ? 9'ha : _GEN_2; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_4 = 6'h4 == instcnt ? 9'h5a : _GEN_3; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_5 = 6'h5 == instcnt ? 9'h12 : _GEN_4; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_6 = 6'h6 == instcnt ? 9'h1a : _GEN_5; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_7 = 6'h7 == instcnt ? 9'h22 : _GEN_6; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_8 = 6'h8 == instcnt ? 9'h2a : _GEN_7; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_9 = 6'h9 == instcnt ? 9'h32 : _GEN_8; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_10 = 6'ha == instcnt ? 9'h3a : _GEN_9; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_11 = 6'hb == instcnt ? 9'h42 : _GEN_10; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_12 = 6'hc == instcnt ? 9'h4 : _GEN_11; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_13 = 6'hd == instcnt ? 9'h4a : _GEN_12; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_14 = 6'he == instcnt ? 9'h82 : _GEN_13; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_15 = 6'hf == instcnt ? 9'hd2 : _GEN_14; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_16 = 6'h10 == instcnt ? 9'h8a : _GEN_15; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_17 = 6'h11 == instcnt ? 9'hda : _GEN_16; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_18 = 6'h12 == instcnt ? 9'h92 : _GEN_17; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_19 = 6'h13 == instcnt ? 9'h9a : _GEN_18; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_20 = 6'h14 == instcnt ? 9'ha2 : _GEN_19; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_21 = 6'h15 == instcnt ? 9'haa : _GEN_20; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_22 = 6'h16 == instcnt ? 9'hb2 : _GEN_21; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_23 = 6'h17 == instcnt ? 9'hba : _GEN_22; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_24 = 6'h18 == instcnt ? 9'hc2 : _GEN_23; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_25 = 6'h19 == instcnt ? 9'h84 : _GEN_24; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_26 = 6'h1a == instcnt ? 9'hca : _GEN_25; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_27 = 6'h1b == instcnt ? 9'h3 : _GEN_26; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_28 = 6'h1c == instcnt ? 9'h13 : _GEN_27; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_29 = 6'h1d == instcnt ? 9'hb : _GEN_28; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_30 = 6'h1e == instcnt ? 9'h1b : _GEN_29; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_31 = 6'h1f == instcnt ? 9'h1c : _GEN_30; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_32 = 6'h20 == instcnt ? 9'h9c : _GEN_31; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_33 = 6'h21 == instcnt ? 9'h152 : _GEN_32; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_34 = 6'h22 == instcnt ? 9'h102 : _GEN_33; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_35 = 6'h23 == instcnt ? 9'h104 : _GEN_34; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_36 = 6'h24 == instcnt ? 9'h14a : _GEN_35; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_37 = 6'h25 == instcnt ? 9'h1d2 : _GEN_36; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_38 = 6'h26 == instcnt ? 9'h182 : _GEN_37; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_39 = 6'h27 == instcnt ? 9'h18a : _GEN_38; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_40 = 6'h28 == instcnt ? 9'h184 : _GEN_39; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_41 = 6'h29 == instcnt ? 9'h1ca : _GEN_40; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_42 = 6'h2a == instcnt ? 9'h103 : _GEN_41; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_43 = 6'h2b == instcnt ? 9'h113 : _GEN_42; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_44 = 6'h2c == instcnt ? 9'h10b : _GEN_43; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_45 = 6'h2d == instcnt ? 9'h11b : _GEN_44; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_46 = 6'h2e == instcnt ? 9'h11c : _GEN_45; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_47 = 6'h2f == instcnt ? 9'h19c : _GEN_46; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_48 = 6'h30 == instcnt ? 9'h62 : _GEN_47; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_49 = 6'h31 == instcnt ? 9'hc : _GEN_48; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_50 = 6'h32 == instcnt ? 9'h14 : _GEN_49; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_51 = 6'h33 == instcnt ? 9'he2 : _GEN_50; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_52 = 6'h34 == instcnt ? 9'h8c : _GEN_51; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_53 = 6'h35 == instcnt ? 9'h94 : _GEN_52; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire [8:0] _GEN_54 = 6'h36 == instcnt ? 9'h1 : _GEN_53; // @[Decodeunit.scala 12:125 Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T = _GEN_54 == 9'h2; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_1 = _GEN_54 == 9'ha; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_2 = _GEN_54 == 9'h12; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_3 = _GEN_54 == 9'h1a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_4 = _GEN_54 == 9'h22; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_5 = _GEN_54 == 9'h2a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_6 = _GEN_54 == 9'h32; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_7 = _GEN_54 == 9'h3a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_8 = _GEN_54 == 9'h42; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_9 = _GEN_54 == 9'h4a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_10 = _GEN_54 == 9'h82; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_11 = _GEN_54 == 9'h8a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_12 = _GEN_54 == 9'h92; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_13 = _GEN_54 == 9'h9a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_14 = _GEN_54 == 9'ha2; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_15 = _GEN_54 == 9'haa; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_16 = _GEN_54 == 9'hb2; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_17 = _GEN_54 == 9'hba; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_18 = _GEN_54 == 9'hc2; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_19 = _GEN_54 == 9'hca; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_20 = _GEN_54 == 9'h102; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_21 = _GEN_54 == 9'h14a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_22 = _GEN_54 == 9'h182; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_23 = _GEN_54 == 9'h18a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_24 = _GEN_54 == 9'h1ca; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_25 = _GEN_54 == 9'h52; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_26 = _GEN_54 == 9'h5a; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_27 = _GEN_54 == 9'h62; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_28 = _GEN_54 == 9'hd2; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_29 = _GEN_54 == 9'hda; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_30 = _GEN_54 == 9'he2; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_31 = _GEN_54 == 9'h152; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_32 = _GEN_54 == 9'h1d2; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_bit_T_33 = _GEN_54 & 9'h11f; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_bit_T_34 = _uop_decoder_bit_T_33 == 9'h13; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_36 = _uop_decoder_bit_T_33 == 9'h113; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_38 = _uop_decoder_bit_T_33 == 9'h1b; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_40 = _uop_decoder_bit_T_33 == 9'h11b; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_41 = _GEN_54 == 9'h4; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_42 = _GEN_54 == 9'h84; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_43 = _GEN_54 == 9'h104; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_44 = _GEN_54 == 9'h184; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_45 = _GEN_54 == 9'h1c; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_46 = _GEN_54 == 9'h9c; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_47 = _GEN_54 == 9'h11c; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_48 = _GEN_54 == 9'h19c; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_49 = _GEN_54 == 9'hc; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_50 = _GEN_54 == 9'h14; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_51 = _GEN_54 == 9'h8c; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_52 = _GEN_54 == 9'h94; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_83 = _uop_decoder_bit_T | _uop_decoder_bit_T_1 | _uop_decoder_bit_T_2 | _uop_decoder_bit_T_3
     | _uop_decoder_bit_T_4 | _uop_decoder_bit_T_5 | _uop_decoder_bit_T_6 | _uop_decoder_bit_T_7 | _uop_decoder_bit_T_8
     | _uop_decoder_bit_T_9 | _uop_decoder_bit_T_10 | _uop_decoder_bit_T_11 | _uop_decoder_bit_T_12 |
    _uop_decoder_bit_T_13 | _uop_decoder_bit_T_14 | _uop_decoder_bit_T_15 | _uop_decoder_bit_T_16 |
    _uop_decoder_bit_T_17 | _uop_decoder_bit_T_18 | _uop_decoder_bit_T_19 | _uop_decoder_bit_T_20 |
    _uop_decoder_bit_T_21 | _uop_decoder_bit_T_22 | _uop_decoder_bit_T_23 | _uop_decoder_bit_T_24 |
    _uop_decoder_bit_T_25 | _uop_decoder_bit_T_26 | _uop_decoder_bit_T_27 | _uop_decoder_bit_T_28 |
    _uop_decoder_bit_T_29 | _uop_decoder_bit_T_30; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_0 = _uop_decoder_bit_T_83 | _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32 | _uop_decoder_bit_T_34 |
    _uop_decoder_bit_T_36 | _uop_decoder_bit_T_38 | _uop_decoder_bit_T_40 | _uop_decoder_bit_T_41 |
    _uop_decoder_bit_T_42 | _uop_decoder_bit_T_43 | _uop_decoder_bit_T_44 | _uop_decoder_bit_T_45 |
    _uop_decoder_bit_T_46 | _uop_decoder_bit_T_47 | _uop_decoder_bit_T_48 | _uop_decoder_bit_T_49 |
    _uop_decoder_bit_T_50 | _uop_decoder_bit_T_51 | _uop_decoder_bit_T_52; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_bit_T_102 = _uop_decoder_bit_T_33 == 9'h3; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_104 = _uop_decoder_bit_T_33 == 9'h103; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_106 = _uop_decoder_bit_T_33 == 9'hb; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_108 = _uop_decoder_bit_T_33 == 9'h10b; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_1 = _uop_decoder_bit_T_102 | _uop_decoder_bit_T_104 | _uop_decoder_bit_T_106 |
    _uop_decoder_bit_T_108; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_bit_T_112 = _GEN_54 & 9'h7; // @[Decodeunit.scala 12:65]
  wire  uop_decoder_2 = _uop_decoder_bit_T_112 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_113 = uop_decoder_2; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_3 = _uop_decoder_bit_T_112 == 9'h1; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_bit_T_115 = uop_decoder_3; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T = _GEN_54 & 9'h8; // @[Decodeunit.scala 12:65]
  wire  uop_decoder_4 = _uop_decoder_T == 9'h8; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_1 = uop_decoder_4; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_2 = _GEN_54 & 9'h9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_3 = _uop_decoder_T_2 == 9'h9; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_4 = _GEN_54 & 9'h48; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_5 = _uop_decoder_T_4 == 9'h48; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_6 = _GEN_54 & 9'h151; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_7 = _uop_decoder_T_6 == 9'h50; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo = _uop_decoder_T_3 | _uop_decoder_T_5 | _uop_decoder_T_7; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_10 = _GEN_54 & 9'h70; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_11 = _uop_decoder_T_10 == 9'h60; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_12 = _GEN_54 & 9'h149; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_13 = _uop_decoder_T_12 == 9'h140; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo = _uop_decoder_T_11 | _uop_decoder_T_13; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_15 = _GEN_54 & 9'h45; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_16 = _uop_decoder_T_15 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_17 = _GEN_54 & 9'h3c; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_18 = _uop_decoder_T_17 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi = _uop_decoder_T_16 | _uop_decoder_T_18; // @[Decodeunit.scala 13:31]
  wire [2:0] uop_decoder_5 = {uop_decoder_hi_hi,uop_decoder_hi_lo,uop_decoder_lo}; // @[Cat.scala 30:58]
  wire  uop_decoder_6 = _uop_decoder_bit_T_38 | _uop_decoder_bit_T_40; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_7 = _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_8 = _uop_decoder_bit_T_34 | _uop_decoder_bit_T_36; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_9 = _uop_decoder_bit_T_9 | _uop_decoder_bit_T_19 | _uop_decoder_bit_T_21 | _uop_decoder_bit_T_24; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_10 = _uop_decoder_bit_T_45 | _uop_decoder_bit_T_46 | _uop_decoder_bit_T_47 | _uop_decoder_bit_T_48; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_20 = _GEN_54 & 9'h100; // @[Decodeunit.scala 12:65]
  wire  uop_decoder_11 = _uop_decoder_T_20 == 9'h100; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_21 = uop_decoder_11; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_12 = _uop_decoder_bit_T_83 | _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32 | _uop_decoder_bit_T_102
     | _uop_decoder_bit_T_104 | _uop_decoder_bit_T_106 | _uop_decoder_bit_T_108 | _uop_decoder_bit_T_34 |
    _uop_decoder_bit_T_36 | _uop_decoder_bit_T_38 | _uop_decoder_bit_T_40 | _uop_decoder_bit_T_41 |
    _uop_decoder_bit_T_42 | _uop_decoder_bit_T_43 | _uop_decoder_bit_T_44 | _uop_decoder_bit_T_45 |
    _uop_decoder_bit_T_46 | _uop_decoder_bit_T_47 | _uop_decoder_bit_T_48 | _uop_decoder_bit_T_49 |
    _uop_decoder_bit_T_50 | _uop_decoder_bit_T_51 | _uop_decoder_bit_T_52; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_22 = _GEN_54 & 9'he9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_23 = _uop_decoder_T_22 == 9'h20; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_24 = _GEN_54 & 9'hf9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_25 = _uop_decoder_T_24 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_26 = _GEN_54 & 9'h1e1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_27 = _uop_decoder_T_26 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_28 = _GEN_54 & 9'he5; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_29 = _uop_decoder_T_28 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_30 = _GEN_54 & 9'h89; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_31 = _uop_decoder_T_30 == 9'h88; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_32 = _GEN_54 & 9'h1b1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_33 = _uop_decoder_T_32 == 9'h90; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_34 = _GEN_54 & 9'he1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_35 = _uop_decoder_T_34 == 9'he0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_36 = _GEN_54 & 9'h109; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_37 = _uop_decoder_T_36 == 9'h109; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_38 = _GEN_54 & 9'h111; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_39 = _uop_decoder_T_38 == 9'h111; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo = _uop_decoder_T_23 | _uop_decoder_T_25 | _uop_decoder_T_27 | _uop_decoder_T_29 |
    _uop_decoder_T_31 | _uop_decoder_T_33 | _uop_decoder_T_35 | _uop_decoder_T_37 | _uop_decoder_T_39; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_48 = _GEN_54 & 9'h102; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_49 = _uop_decoder_T_48 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_50 = _GEN_54 & 9'h101; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_51 = _uop_decoder_T_50 == 9'h1; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_52 = _GEN_54 & 9'h118; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_53 = _uop_decoder_T_52 == 9'h8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_54 = _GEN_54 & 9'h98; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_55 = _uop_decoder_T_54 == 9'h10; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_56 = _GEN_54 & 9'h11; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_57 = _uop_decoder_T_56 == 9'h11; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_58 = _GEN_54 & 9'h160; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_59 = _uop_decoder_T_58 == 9'h60; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_60 = _GEN_54 & 9'h190; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_61 = _uop_decoder_T_60 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_62 = _GEN_54 & 9'h92; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_63 = _uop_decoder_T_62 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_64 = _GEN_54 & 9'h170; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_65 = _uop_decoder_T_64 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_66 = _GEN_54 & 9'h138; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_67 = _uop_decoder_T_66 == 9'h10; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_lo = _uop_decoder_T_49 | _uop_decoder_T_51 | _uop_decoder_T_53 | _uop_decoder_T_3 |
    _uop_decoder_T_55 | _uop_decoder_T_57 | _uop_decoder_T_59 | _uop_decoder_T_61 | _uop_decoder_T_63 |
    _uop_decoder_T_65 | _uop_decoder_T_67; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_78 = _GEN_54 & 9'h131; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_79 = _uop_decoder_T_78 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_80 = _GEN_54 & 9'h129; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_81 = _uop_decoder_T_80 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_82 = _GEN_54 & 9'h39; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_83 = _uop_decoder_T_82 == 9'h38; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_84 = _GEN_54 & 9'h141; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_85 = _uop_decoder_T_84 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_86 = _GEN_54 & 9'h49; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_87 = _uop_decoder_T_86 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_88 = _GEN_54 & 9'h119; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_89 = _uop_decoder_T_88 == 9'h101; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_90 = _GEN_54 & 9'h99; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_91 = _uop_decoder_T_90 == 9'h90; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_hi = _uop_decoder_T_79 | _uop_decoder_T_81 | _uop_decoder_T_49 | _uop_decoder_T_83 |
    _uop_decoder_T_85 | _uop_decoder_T_87 | _uop_decoder_T_89 | _uop_decoder_T_91; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_99 = _GEN_54 & 9'h19; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_100 = _uop_decoder_T_99 == 9'h1; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_101 = _GEN_54 & 9'hd9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_102 = _uop_decoder_T_101 == 9'h50; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_103 = _GEN_54 & 9'h19a; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_104 = _uop_decoder_T_103 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_105 = _GEN_54 & 9'hdd; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_106 = _uop_decoder_T_105 == 9'h98; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_108 = _uop_decoder_T_34 == 9'ha0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_109 = _GEN_54 & 9'hf8; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_110 = _uop_decoder_T_109 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_1 = _uop_decoder_T_100 | _uop_decoder_T_102 | _uop_decoder_T_104 | _uop_decoder_T_106 |
    _uop_decoder_T_108 | _uop_decoder_T_110; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_116 = _GEN_54 & 9'h11a; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_117 = _uop_decoder_T_116 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_118 = _GEN_54 & 9'h5d; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_119 = _uop_decoder_T_118 == 9'h18; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_120 = _GEN_54 & 9'h61; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_121 = _uop_decoder_T_120 == 9'h20; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_122 = _GEN_54 & 9'h79; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_123 = _uop_decoder_T_122 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_124 = _GEN_54 & 9'h1e9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_125 = _uop_decoder_T_124 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_lo = _uop_decoder_T_117 | _uop_decoder_T_119 | _uop_decoder_T_121 | _uop_decoder_T_123 |
    _uop_decoder_T_125; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_130 = _GEN_54 & 9'h112; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_131 = _uop_decoder_T_130 == 9'h100; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_132 = _GEN_54 & 9'h159; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_133 = _uop_decoder_T_132 == 9'h108; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_hi = _uop_decoder_T_131 | _uop_decoder_T_133; // @[Decodeunit.scala 13:31]
  wire [5:0] uop_decoder_15 = {uop_decoder_hi_hi_hi,uop_decoder_hi_hi_lo,uop_decoder_hi_lo_1,uop_decoder_lo_hi_hi,
    uop_decoder_lo_hi_lo,uop_decoder_lo_lo}; // @[Cat.scala 30:58]
  wire  uop_decoder_16 = _uop_decoder_bit_T_83 | _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32 | _uop_decoder_bit_T_38
     | _uop_decoder_bit_T_40; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_135 = _GEN_54 & 9'h41; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_136 = _uop_decoder_T_135 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_137 = _GEN_54 & 9'h38; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_138 = _uop_decoder_T_137 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_17 = _uop_decoder_T_136 | _uop_decoder_T_138; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_140 = _GEN_54 & 9'hc9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_141 = _uop_decoder_T_140 == 9'h8; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_143 = _uop_decoder_T_90 == 9'h18; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_144 = _GEN_54 & 9'hf0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_145 = _uop_decoder_T_144 == 9'h60; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_146 = _GEN_54 & 9'hc8; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_147 = _uop_decoder_T_146 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_149 = _uop_decoder_T_144 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_150 = _GEN_54 & 9'h110; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_151 = _uop_decoder_T_150 == 9'h110; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo_1 = _uop_decoder_T_141 | _uop_decoder_T_143 | _uop_decoder_T_145 | _uop_decoder_T_147 |
    _uop_decoder_T_149 | _uop_decoder_T_151; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_158 = _uop_decoder_T_60 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_159 = _GEN_54 & 9'h158; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_160 = _uop_decoder_T_159 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_162 = _uop_decoder_T_64 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_163 = _GEN_54 & 9'h1c9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_164 = _uop_decoder_T_163 == 9'h48; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_166 = _uop_decoder_T_101 == 9'h98; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_168 = _uop_decoder_T_159 == 9'h108; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_169 = _GEN_54 & 9'h1c8; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_170 = _uop_decoder_T_169 == 9'h140; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_lo_1 = _uop_decoder_T_158 | _uop_decoder_T_160 | _uop_decoder_T_162 | _uop_decoder_T_164 |
    _uop_decoder_T_166 | _uop_decoder_T_168 | _uop_decoder_T_170; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_177 = _GEN_54 & 9'h1f0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_178 = _uop_decoder_T_177 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_180 = _uop_decoder_T_66 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_181 = _GEN_54 & 9'h31; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_182 = _uop_decoder_T_181 == 9'h30; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_183 = _GEN_54 & 9'hd8; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_184 = _uop_decoder_T_183 == 9'h40; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_186 = _uop_decoder_T_101 == 9'h58; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_187 = _GEN_54 & 9'ha9; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_188 = _uop_decoder_T_187 == 9'ha8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_189 = _GEN_54 & 9'h150; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_190 = _uop_decoder_T_189 == 9'h140; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_191 = _GEN_54 & 9'h148; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_192 = _uop_decoder_T_191 == 9'h140; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_hi_1 = _uop_decoder_T_178 | _uop_decoder_T_180 | _uop_decoder_T_182 | _uop_decoder_T_184 |
    _uop_decoder_T_186 | _uop_decoder_T_188 | _uop_decoder_T_190 | _uop_decoder_T_192; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_200 = _GEN_54 & 9'h1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_201 = _uop_decoder_T_200 == 9'h1; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_202 = _GEN_54 & 9'hd0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_203 = _uop_decoder_T_202 == 9'h90; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_204 = _GEN_54 & 9'he0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_205 = _uop_decoder_T_204 == 9'ha0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_206 = _GEN_54 & 9'h188; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_207 = _uop_decoder_T_206 == 9'h88; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_2 = _uop_decoder_T_178 | _uop_decoder_T_201 | _uop_decoder_T_5 | _uop_decoder_T_203 |
    _uop_decoder_T_205 | _uop_decoder_T_149 | _uop_decoder_T_207; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_214 = _GEN_54 & 9'h51; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_215 = _uop_decoder_T_214 == 9'h10; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_216 = _GEN_54 & 9'h78; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_217 = _uop_decoder_T_216 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_218 = _GEN_54 & 9'h1c1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_219 = _uop_decoder_T_218 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_221 = _uop_decoder_T_90 == 9'h98; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_lo_1 = _uop_decoder_T_215 | _uop_decoder_T_121 | _uop_decoder_T_217 | _uop_decoder_T_219 |
    _uop_decoder_T_221 | _uop_decoder_T_170; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_228 = _uop_decoder_T_159 == 9'h50; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_230 = _uop_decoder_T_189 == 9'h100; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_hi_1 = _uop_decoder_T_228 | _uop_decoder_T_230; // @[Decodeunit.scala 13:31]
  wire [5:0] uop_decoder_19 = {uop_decoder_hi_hi_hi_1,uop_decoder_hi_hi_lo_1,uop_decoder_hi_lo_2,uop_decoder_lo_hi_hi_1,
    uop_decoder_lo_hi_lo_1,uop_decoder_lo_lo_1}; // @[Cat.scala 30:58]
  wire  uop_decoder_20 = _uop_decoder_bit_T | _uop_decoder_bit_T_1 | _uop_decoder_bit_T_2 | _uop_decoder_bit_T_3 |
    _uop_decoder_bit_T_4 | _uop_decoder_bit_T_5 | _uop_decoder_bit_T_6 | _uop_decoder_bit_T_7 | _uop_decoder_bit_T_8 |
    _uop_decoder_bit_T_10 | _uop_decoder_bit_T_11 | _uop_decoder_bit_T_12 | _uop_decoder_bit_T_13 |
    _uop_decoder_bit_T_14 | _uop_decoder_bit_T_15 | _uop_decoder_bit_T_16 | _uop_decoder_bit_T_17 |
    _uop_decoder_bit_T_18 | _uop_decoder_bit_T_20 | _uop_decoder_bit_T_22 | _uop_decoder_bit_T_23 |
    _uop_decoder_bit_T_27 | _uop_decoder_bit_T_30 | _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32 |
    _uop_decoder_bit_T_38 | _uop_decoder_bit_T_40; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_232 = _GEN_54 & 9'h30; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_233 = _uop_decoder_T_232 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_21 = _uop_decoder_T_136 | _uop_decoder_T_233; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_236 = _uop_decoder_T_30 == 9'h8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_237 = _GEN_54 & 9'h88; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_238 = _uop_decoder_T_237 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_240 = _uop_decoder_T_52 == 9'h118; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo_2 = _uop_decoder_T_236 | _uop_decoder_T_11 | _uop_decoder_T_238 | _uop_decoder_T_240; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_244 = _GEN_54 & 9'h1d0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_245 = _uop_decoder_T_244 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_247 = _uop_decoder_T_204 == 9'h40; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_249 = _uop_decoder_T_54 == 9'h98; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_250 = _GEN_54 & 9'h108; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_251 = _uop_decoder_T_250 == 9'h108; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_lo_2 = _uop_decoder_T_245 | _uop_decoder_T_160 | _uop_decoder_T_180 | _uop_decoder_T_201 |
    _uop_decoder_T_247 | _uop_decoder_T_249 | _uop_decoder_T_251; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_258 = _GEN_54 & 9'h1b0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_259 = _uop_decoder_T_258 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_260 = _GEN_54 & 9'h68; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_261 = _uop_decoder_T_260 == 9'h40; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_hi_2 = _uop_decoder_T_259 | _uop_decoder_T_180 | _uop_decoder_T_182 | _uop_decoder_T_261 |
    _uop_decoder_T_188; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_266 = _GEN_54 & 9'h191; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_267 = _uop_decoder_T_266 == 9'h90; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_269 = _uop_decoder_T_66 == 9'h8; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_3 = _uop_decoder_T_178 | _uop_decoder_T_267 | _uop_decoder_T_108 | _uop_decoder_T_149 |
    _uop_decoder_T_170 | _uop_decoder_T_269; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_276 = _uop_decoder_T_56 == 9'h10; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_278 = _uop_decoder_T_10 == 9'h40; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_lo_2 = _uop_decoder_T_276 | _uop_decoder_T_121 | _uop_decoder_T_278 | _uop_decoder_T_219; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_hi_hi_hi_2 = _uop_decoder_T_150 == 9'h100; // @[Decodeunit.scala 12:125]
  wire [5:0] uop_decoder_23 = {uop_decoder_hi_hi_hi_2,uop_decoder_hi_hi_lo_2,uop_decoder_hi_lo_3,uop_decoder_lo_hi_hi_2,
    uop_decoder_lo_hi_lo_2,uop_decoder_lo_lo_2}; // @[Cat.scala 30:58]
  wire  uop_decoder_24 = _uop_decoder_bit_T | _uop_decoder_bit_T_1 | _uop_decoder_bit_T_2 | _uop_decoder_bit_T_3 |
    _uop_decoder_bit_T_4 | _uop_decoder_bit_T_5 | _uop_decoder_bit_T_6 | _uop_decoder_bit_T_7 | _uop_decoder_bit_T_8 |
    _uop_decoder_bit_T_10 | _uop_decoder_bit_T_11 | _uop_decoder_bit_T_12 | _uop_decoder_bit_T_13 |
    _uop_decoder_bit_T_14 | _uop_decoder_bit_T_15 | _uop_decoder_bit_T_16 | _uop_decoder_bit_T_17 |
    _uop_decoder_bit_T_18 | _uop_decoder_bit_T_20 | _uop_decoder_bit_T_22 | _uop_decoder_bit_T_23 |
    _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_285 = _uop_decoder_T_20 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_286 = _GEN_54 & 9'h40; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_287 = _uop_decoder_T_286 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_25 = _uop_decoder_T_285 | _uop_decoder_T_287; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_290 = _uop_decoder_T_237 == 9'h8; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_292 = _uop_decoder_T_206 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_293 = _GEN_54 & 9'h1c0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_294 = _uop_decoder_T_293 == 9'h140; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo_3 = _uop_decoder_T_290 | _uop_decoder_T_292 | _uop_decoder_T_147 | _uop_decoder_T_294; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_299 = _uop_decoder_T_52 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_301 = _uop_decoder_T_286 == 9'h40; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_lo_3 = _uop_decoder_T_158 | _uop_decoder_T_299 | _uop_decoder_T_301 | _uop_decoder_T_249 |
    _uop_decoder_T_251; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_307 = _uop_decoder_T_232 == 9'h30; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_308 = _GEN_54 & 9'ha8; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_309 = _uop_decoder_T_308 == 9'ha8; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_hi_3 = _uop_decoder_T_259 | _uop_decoder_T_180 | _uop_decoder_T_307 | _uop_decoder_T_301 |
    _uop_decoder_T_309; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_315 = _uop_decoder_T_60 == 9'h90; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_316 = _GEN_54 & 9'ha0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_317 = _uop_decoder_T_316 == 9'ha0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_319 = _uop_decoder_T_293 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_4 = _uop_decoder_T_178 | _uop_decoder_T_315 | _uop_decoder_T_317 | _uop_decoder_T_319 |
    _uop_decoder_T_294 | _uop_decoder_T_207; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_325 = _GEN_54 & 9'h10; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_326 = _uop_decoder_T_325 == 9'h10; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_327 = _GEN_54 & 9'h20; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_328 = _uop_decoder_T_327 == 9'h20; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_329 = _GEN_54 & 9'h180; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_330 = _uop_decoder_T_329 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_lo_3 = _uop_decoder_T_326 | _uop_decoder_T_328 | _uop_decoder_T_301 | _uop_decoder_T_330; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_334 = _GEN_54 & 9'h140; // @[Decodeunit.scala 12:65]
  wire  uop_decoder_hi_hi_hi_3 = _uop_decoder_T_334 == 9'h100; // @[Decodeunit.scala 12:125]
  wire [5:0] uop_decoder_27 = {uop_decoder_hi_hi_hi_3,uop_decoder_hi_hi_lo_3,uop_decoder_hi_lo_4,uop_decoder_lo_hi_hi_3,
    uop_decoder_lo_hi_lo_3,uop_decoder_lo_lo_3}; // @[Cat.scala 30:58]
  wire  _uop_decoder_T_337 = 1'h1; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo_4 = _uop_decoder_T_290 | _uop_decoder_T_238; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_lo_hi_lo_4 = _uop_decoder_T_158 | _uop_decoder_T_299 | _uop_decoder_T_249 | _uop_decoder_T_251; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_lo_hi_hi_4 = _uop_decoder_T_259 | _uop_decoder_T_180 | _uop_decoder_T_307 | _uop_decoder_T_309; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_345 = _GEN_54 & 9'h90; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_346 = _uop_decoder_T_345 == 9'h90; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_347 = _GEN_54 & 9'hc0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_348 = _uop_decoder_T_347 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_5 = _uop_decoder_T_178 | _uop_decoder_T_346 | _uop_decoder_T_317 | _uop_decoder_T_348 |
    _uop_decoder_T_207; // @[Decodeunit.scala 13:31]
  wire [5:0] uop_decoder_31 = {uop_decoder_11,uop_decoder_hi_hi_lo_3,uop_decoder_hi_lo_5,uop_decoder_lo_hi_hi_4,
    uop_decoder_lo_hi_lo_4,uop_decoder_lo_lo_4}; // @[Cat.scala 30:58]
  wire  uop_decoder_32 = _uop_decoder_bit_T_83 | _uop_decoder_bit_T_31 | _uop_decoder_bit_T_32 | _uop_decoder_bit_T_102
     | _uop_decoder_bit_T_104 | _uop_decoder_bit_T_34 | _uop_decoder_bit_T_36 | _uop_decoder_bit_T_38 |
    _uop_decoder_bit_T_40 | _uop_decoder_bit_T_41 | _uop_decoder_bit_T_42 | _uop_decoder_bit_T_43 |
    _uop_decoder_bit_T_44 | _uop_decoder_bit_T_45 | _uop_decoder_bit_T_46 | _uop_decoder_bit_T_47 |
    _uop_decoder_bit_T_48 | _uop_decoder_bit_T_49 | _uop_decoder_bit_T_50 | _uop_decoder_bit_T_51 |
    _uop_decoder_bit_T_52; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_356 = _GEN_54 & 9'h5; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_357 = _uop_decoder_T_356 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_358 = _GEN_54 & 9'hc; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_359 = _uop_decoder_T_358 == 9'h8; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_33 = _uop_decoder_T_357 | _uop_decoder_T_359; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_361 = _GEN_54 & 9'h14; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_362 = _uop_decoder_T_361 == 9'h10; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_364 = _uop_decoder_T_56 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_365 = _GEN_54 & 9'ha; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_366 = _uop_decoder_T_365 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_34 = _uop_decoder_T_362 | _uop_decoder_T_364 | _uop_decoder_T_366; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_370 = _uop_decoder_T_62 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_372 = _uop_decoder_T_36 == 9'h1; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_374 = _uop_decoder_T_56 == 9'h1; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_375 = _GEN_54 & 9'hcd; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_376 = _uop_decoder_T_375 == 9'h8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_377 = _GEN_54 & 9'h1a; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_378 = _uop_decoder_T_377 == 9'h8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_379 = _GEN_54 & 9'h1cc; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_380 = _uop_decoder_T_379 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_382 = _uop_decoder_T_140 == 9'hc8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_383 = _GEN_54 & 9'hbc; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_384 = _uop_decoder_T_383 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo_5 = _uop_decoder_T_370 | _uop_decoder_T_372 | _uop_decoder_T_374 | _uop_decoder_T_376 |
    _uop_decoder_T_378 | _uop_decoder_T_102 | _uop_decoder_T_145 | _uop_decoder_T_380 | _uop_decoder_T_382 |
    _uop_decoder_T_240 | _uop_decoder_T_384; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_395 = _GEN_54 & 9'h15c; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_396 = _uop_decoder_T_395 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_398 = _uop_decoder_T_38 == 9'h1; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_399 = _GEN_54 & 9'h169; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_400 = _uop_decoder_T_399 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_401 = _GEN_54 & 9'h9d; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_402 = _uop_decoder_T_401 == 9'h98; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_404 = _uop_decoder_T_22 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_406 = _uop_decoder_T_88 == 9'h111; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_407 = _GEN_54 & 9'h192; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_408 = _uop_decoder_T_407 == 9'h180; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_lo_5 = _uop_decoder_T_245 | _uop_decoder_T_396 | _uop_decoder_T_398 | _uop_decoder_T_378 |
    _uop_decoder_T_400 | _uop_decoder_T_402 | _uop_decoder_T_404 | _uop_decoder_T_168 | _uop_decoder_T_406 |
    _uop_decoder_T_408 | _uop_decoder_T_162; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_419 = _GEN_54 & 9'h1f5; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_420 = _uop_decoder_T_419 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_421 = _GEN_54 & 9'h13d; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_422 = _uop_decoder_T_421 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_424 = _uop_decoder_T_101 == 9'h40; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_425 = _GEN_54 & 9'h59; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_426 = _uop_decoder_T_425 == 9'h58; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_428 = _uop_decoder_T_38 == 9'h101; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_429 = _GEN_54 & 9'h1d1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_430 = _uop_decoder_T_429 == 9'hd0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_hi_5 = _uop_decoder_T_420 | _uop_decoder_T_422 | _uop_decoder_T_378 | _uop_decoder_T_182 |
    _uop_decoder_T_424 | _uop_decoder_T_426 | _uop_decoder_T_63 | _uop_decoder_T_188 | _uop_decoder_T_131 |
    _uop_decoder_T_428 | _uop_decoder_T_190 | _uop_decoder_T_430; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_442 = _GEN_54 & 9'h12; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_443 = _uop_decoder_T_442 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_445 = _uop_decoder_T_365 == 9'h8; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_446 = _GEN_54 & 9'hd5; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_447 = _uop_decoder_T_446 == 9'h90; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_449 = _uop_decoder_T_202 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_451 = _uop_decoder_T_84 == 9'h140; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_452 = _GEN_54 & 9'hb0; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_453 = _uop_decoder_T_452 == 9'ha0; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_6 = _uop_decoder_T_178 | _uop_decoder_T_443 | _uop_decoder_T_374 | _uop_decoder_T_445 |
    _uop_decoder_T_3 | _uop_decoder_T_447 | _uop_decoder_T_449 | _uop_decoder_T_451 | _uop_decoder_T_269 |
    _uop_decoder_T_453; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_463 = _GEN_54 & 9'h58; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_464 = _uop_decoder_T_463 == 9'h10; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_465 = _GEN_54 & 9'h55; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_466 = _uop_decoder_T_465 == 9'h10; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_468 = _uop_decoder_T_99 == 9'h11; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_469 = _GEN_54 & 9'h1c5; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_470 = _uop_decoder_T_469 == 9'h80; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_lo_5 = _uop_decoder_T_464 | _uop_decoder_T_466 | _uop_decoder_T_468 | _uop_decoder_T_121 |
    _uop_decoder_T_123 | _uop_decoder_T_470; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_477 = _uop_decoder_T_214 == 9'h50; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_479 = _uop_decoder_T_120 == 9'h60; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_481 = _uop_decoder_T_6 == 9'h100; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_hi_hi_5 = _uop_decoder_T_443 | _uop_decoder_T_366 | _uop_decoder_T_468 | _uop_decoder_T_477 |
    _uop_decoder_T_479 | _uop_decoder_T_481; // @[Decodeunit.scala 13:31]
  wire [5:0] uop_decoder_35 = {uop_decoder_hi_hi_hi_5,uop_decoder_hi_hi_lo_5,uop_decoder_hi_lo_6,uop_decoder_lo_hi_hi_5,
    uop_decoder_lo_hi_lo_5,uop_decoder_lo_lo_5}; // @[Cat.scala 30:58]
  wire  _uop_decoder_T_488 = _uop_decoder_T_30 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_489 = _GEN_54 & 9'h82; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_490 = _uop_decoder_T_489 == 9'h80; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_491 = _GEN_54 & 9'hc1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_492 = _uop_decoder_T_491 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_494 = _uop_decoder_T_50 == 9'h101; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_lo_6 = _uop_decoder_T_376 | _uop_decoder_T_488 | _uop_decoder_T_490 | _uop_decoder_T_492 |
    _uop_decoder_T_494; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_500 = _uop_decoder_T_2 == 9'h1; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_501 = _GEN_54 & 9'h199; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_502 = _uop_decoder_T_501 == 9'h98; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_lo_6 = _uop_decoder_T_158 | _uop_decoder_T_299 | _uop_decoder_T_49 | _uop_decoder_T_374 |
    _uop_decoder_T_500 | _uop_decoder_T_85 | _uop_decoder_T_502 | _uop_decoder_T_168; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_510 = _GEN_54 & 9'h1f1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_511 = _uop_decoder_T_510 == 9'h0; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_512 = _GEN_54 & 9'h139; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_513 = _uop_decoder_T_512 == 9'h0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_515 = _uop_decoder_T_12 == 9'h40; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_517 = _uop_decoder_T_6 == 9'h140; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_lo_hi_hi_6 = _uop_decoder_T_511 | _uop_decoder_T_513 | _uop_decoder_T_49 | _uop_decoder_T_182 |
    _uop_decoder_T_515 | _uop_decoder_T_7 | _uop_decoder_T_188 | _uop_decoder_T_517; // @[Decodeunit.scala 13:31]
  wire  _uop_decoder_T_526 = _uop_decoder_T_99 == 9'h19; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_528 = _uop_decoder_T_425 == 9'h48; // @[Decodeunit.scala 12:125]
  wire [8:0] _uop_decoder_T_529 = _GEN_54 & 9'hf1; // @[Decodeunit.scala 12:65]
  wire  _uop_decoder_T_530 = _uop_decoder_T_529 == 9'hc0; // @[Decodeunit.scala 12:125]
  wire  _uop_decoder_T_532 = _uop_decoder_T_421 == 9'h8; // @[Decodeunit.scala 12:125]
  wire  uop_decoder_hi_lo_7 = _uop_decoder_T_420 | _uop_decoder_T_526 | _uop_decoder_T_528 | _uop_decoder_T_447 |
    _uop_decoder_T_108 | _uop_decoder_T_530 | _uop_decoder_T_532; // @[Decodeunit.scala 13:31]
  wire  uop_decoder_hi_hi_lo_6 = _uop_decoder_T_466 | _uop_decoder_T_121 | _uop_decoder_T_123 | _uop_decoder_T_470; // @[Decodeunit.scala 13:31]
  wire [8:0] _uop_decoder_T_542 = _GEN_54 & 9'h145; // @[Decodeunit.scala 12:65]
  wire  uop_decoder_hi_hi_hi_6 = _uop_decoder_T_542 == 9'h100; // @[Decodeunit.scala 12:125]
  wire [5:0] uop_decoder_37 = {uop_decoder_hi_hi_hi_6,uop_decoder_hi_hi_lo_6,uop_decoder_hi_lo_7,uop_decoder_lo_hi_hi_6,
    uop_decoder_lo_hi_lo_6,uop_decoder_lo_lo_6}; // @[Cat.scala 30:58]
  wire  uop_srcreq_0_iscoef = 1'h0; // @[dspdecode.scala 76:17 decode.scala 116:42]
  wire  uop_srcreq_0_valid = uop_decoder_12; // @[Decodeunit.scala 13:31]
  wire  vld = uop_srcreq_0_valid & ~uop_srcreq_0_iscoef; // @[dspdecode.scala 81:35]
  wire [5:0] uop_srcreq_0_idx = uop_decoder_15; // @[Cat.scala 30:58]
  wire  idx__0 = vld & io_wd_check_0_valid & uop_srcreq_0_idx == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  wire  idx__1 = vld & io_wd_check_1_valid & uop_srcreq_0_idx == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  wire  idx__2 = vld & io_wd_check_2_valid & uop_srcreq_0_idx == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  wire  idx__3 = vld & io_wd_check_3_valid & uop_srcreq_0_idx == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  wire  idx__4 = vld & io_wd_check_4_valid & uop_srcreq_0_idx == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  wire  idx__5 = vld & io_wd_check_5_valid & uop_srcreq_0_idx == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  wire  _T_2 = idx__0; // @[dspdecode.scala 44:43]
  wire  _T_5 = idx__1; // @[dspdecode.scala 44:43]
  wire  _T_8 = idx__2; // @[dspdecode.scala 44:43]
  wire  _T_11 = idx__3; // @[dspdecode.scala 44:43]
  wire  _T_14 = idx__4; // @[dspdecode.scala 44:43]
  wire  _T_17 = idx__5; // @[dspdecode.scala 44:43]
  wire  busy = idx__0 | idx__1 | idx__2 | idx__3 | idx__4 | idx__5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_1_iscoef = 1'h0; // @[dspdecode.scala 76:17 decode.scala 116:42]
  wire  uop_srcreq_1_valid = uop_decoder_16; // @[Decodeunit.scala 13:31]
  wire  vld_1 = uop_srcreq_1_valid & ~uop_srcreq_0_iscoef; // @[dspdecode.scala 81:35]
  wire [5:0] uop_srcreq_1_idx = uop_decoder_19; // @[Cat.scala 30:58]
  wire  idx_1_0 = vld_1 & io_wd_check_0_valid & uop_srcreq_1_idx == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  wire  idx_1_1 = vld_1 & io_wd_check_1_valid & uop_srcreq_1_idx == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  wire  idx_1_2 = vld_1 & io_wd_check_2_valid & uop_srcreq_1_idx == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  wire  idx_1_3 = vld_1 & io_wd_check_3_valid & uop_srcreq_1_idx == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  wire  idx_1_4 = vld_1 & io_wd_check_4_valid & uop_srcreq_1_idx == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  wire  idx_1_5 = vld_1 & io_wd_check_5_valid & uop_srcreq_1_idx == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  wire  _T_20 = idx_1_0; // @[dspdecode.scala 44:43]
  wire  _T_23 = idx_1_1; // @[dspdecode.scala 44:43]
  wire  _T_26 = idx_1_2; // @[dspdecode.scala 44:43]
  wire  _T_29 = idx_1_3; // @[dspdecode.scala 44:43]
  wire  _T_32 = idx_1_4; // @[dspdecode.scala 44:43]
  wire  _T_35 = idx_1_5; // @[dspdecode.scala 44:43]
  wire  busy_1 = idx_1_0 | idx_1_1 | idx_1_2 | idx_1_3 | idx_1_4 | idx_1_5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_2_iscoef = 1'h0; // @[dspdecode.scala 76:17 decode.scala 116:42]
  wire  uop_srcreq_2_valid = uop_decoder_20; // @[Decodeunit.scala 13:31]
  wire  vld_2 = uop_srcreq_2_valid & ~uop_srcreq_0_iscoef; // @[dspdecode.scala 81:35]
  wire [5:0] uop_srcreq_2_idx = uop_decoder_23; // @[Cat.scala 30:58]
  wire  idx_2_0 = vld_2 & io_wd_check_0_valid & uop_srcreq_2_idx == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  wire  idx_2_1 = vld_2 & io_wd_check_1_valid & uop_srcreq_2_idx == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  wire  idx_2_2 = vld_2 & io_wd_check_2_valid & uop_srcreq_2_idx == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  wire  idx_2_3 = vld_2 & io_wd_check_3_valid & uop_srcreq_2_idx == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  wire  idx_2_4 = vld_2 & io_wd_check_4_valid & uop_srcreq_2_idx == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  wire  idx_2_5 = vld_2 & io_wd_check_5_valid & uop_srcreq_2_idx == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  wire  _T_38 = idx_2_0; // @[dspdecode.scala 44:43]
  wire  _T_41 = idx_2_1; // @[dspdecode.scala 44:43]
  wire  _T_44 = idx_2_2; // @[dspdecode.scala 44:43]
  wire  _T_47 = idx_2_3; // @[dspdecode.scala 44:43]
  wire  _T_50 = idx_2_4; // @[dspdecode.scala 44:43]
  wire  _T_53 = idx_2_5; // @[dspdecode.scala 44:43]
  wire  busy_2 = idx_2_0 | idx_2_1 | idx_2_2 | idx_2_3 | idx_2_4 | idx_2_5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_3_iscoef = 1'h0; // @[dspdecode.scala 76:17 decode.scala 116:42]
  wire  uop_srcreq_3_valid = uop_decoder_24; // @[Decodeunit.scala 13:31]
  wire  vld_3 = uop_srcreq_3_valid & ~uop_srcreq_0_iscoef; // @[dspdecode.scala 81:35]
  wire [5:0] uop_srcreq_3_idx = uop_decoder_27; // @[Cat.scala 30:58]
  wire  idx_3_0 = vld_3 & io_wd_check_0_valid & uop_srcreq_3_idx == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  wire  idx_3_1 = vld_3 & io_wd_check_1_valid & uop_srcreq_3_idx == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  wire  idx_3_2 = vld_3 & io_wd_check_2_valid & uop_srcreq_3_idx == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  wire  idx_3_3 = vld_3 & io_wd_check_3_valid & uop_srcreq_3_idx == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  wire  idx_3_4 = vld_3 & io_wd_check_4_valid & uop_srcreq_3_idx == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  wire  idx_3_5 = vld_3 & io_wd_check_5_valid & uop_srcreq_3_idx == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  wire  _T_56 = idx_3_0; // @[dspdecode.scala 44:43]
  wire  _T_59 = idx_3_1; // @[dspdecode.scala 44:43]
  wire  _T_62 = idx_3_2; // @[dspdecode.scala 44:43]
  wire  _T_65 = idx_3_3; // @[dspdecode.scala 44:43]
  wire  _T_68 = idx_3_4; // @[dspdecode.scala 44:43]
  wire  _T_71 = idx_3_5; // @[dspdecode.scala 44:43]
  wire  busy_3 = idx_3_0 | idx_3_1 | idx_3_2 | idx_3_3 | idx_3_4 | idx_3_5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_4_iscoef = 1'h0; // @[dspdecode.scala 76:17 decode.scala 116:42]
  wire  uop_srcreq_4_valid = _uop_decoder_bit_T | _uop_decoder_bit_T_1 | _uop_decoder_bit_T_2 | _uop_decoder_bit_T_3 |
    _uop_decoder_bit_T_4 | _uop_decoder_bit_T_5 | _uop_decoder_bit_T_6 | _uop_decoder_bit_T_7 | _uop_decoder_bit_T_8 |
    _uop_decoder_bit_T_10 | _uop_decoder_bit_T_11 | _uop_decoder_bit_T_12 | _uop_decoder_bit_T_13 |
    _uop_decoder_bit_T_14 | _uop_decoder_bit_T_15 | _uop_decoder_bit_T_16 | _uop_decoder_bit_T_17 |
    _uop_decoder_bit_T_18 | _uop_decoder_bit_T_20 | _uop_decoder_bit_T_22 | _uop_decoder_bit_T_23; // @[Decodeunit.scala 13:31]
  wire  vld_4 = uop_srcreq_4_valid & ~uop_srcreq_0_iscoef; // @[dspdecode.scala 81:35]
  wire [5:0] uop_srcreq_4_idx = uop_decoder_31; // @[Cat.scala 30:58]
  wire  idx_4_0 = vld_4 & io_wd_check_0_valid & uop_srcreq_4_idx == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  wire  idx_4_1 = vld_4 & io_wd_check_1_valid & uop_srcreq_4_idx == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  wire  idx_4_2 = vld_4 & io_wd_check_2_valid & uop_srcreq_4_idx == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  wire  idx_4_3 = vld_4 & io_wd_check_3_valid & uop_srcreq_4_idx == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  wire  idx_4_4 = vld_4 & io_wd_check_4_valid & uop_srcreq_4_idx == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  wire  idx_4_5 = vld_4 & io_wd_check_5_valid & uop_srcreq_4_idx == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  wire  _T_74 = idx_4_0; // @[dspdecode.scala 44:43]
  wire  _T_77 = idx_4_1; // @[dspdecode.scala 44:43]
  wire  _T_80 = idx_4_2; // @[dspdecode.scala 44:43]
  wire  _T_83 = idx_4_3; // @[dspdecode.scala 44:43]
  wire  _T_86 = idx_4_4; // @[dspdecode.scala 44:43]
  wire  _T_89 = idx_4_5; // @[dspdecode.scala 44:43]
  wire  busy_4 = idx_4_0 | idx_4_1 | idx_4_2 | idx_4_3 | idx_4_4 | idx_4_5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_5_iscoef = uop_decoder_34; // @[Decodeunit.scala 13:31]
  wire  uop_srcreq_5_valid = uop_decoder_32; // @[Decodeunit.scala 13:31]
  wire  vld_5 = uop_srcreq_5_valid & ~uop_srcreq_5_iscoef; // @[dspdecode.scala 81:35]
  wire [5:0] uop_srcreq_5_idx = uop_decoder_35; // @[Cat.scala 30:58]
  wire  idx_5_0 = vld_5 & io_wd_check_0_valid & uop_srcreq_5_idx == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  wire  idx_5_1 = vld_5 & io_wd_check_1_valid & uop_srcreq_5_idx == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  wire  idx_5_2 = vld_5 & io_wd_check_2_valid & uop_srcreq_5_idx == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  wire  idx_5_3 = vld_5 & io_wd_check_3_valid & uop_srcreq_5_idx == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  wire  idx_5_4 = vld_5 & io_wd_check_4_valid & uop_srcreq_5_idx == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  wire  idx_5_5 = vld_5 & io_wd_check_5_valid & uop_srcreq_5_idx == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  wire  _T_92 = idx_5_0; // @[dspdecode.scala 44:43]
  wire  _T_95 = idx_5_1; // @[dspdecode.scala 44:43]
  wire  _T_98 = idx_5_2; // @[dspdecode.scala 44:43]
  wire  _T_101 = idx_5_3; // @[dspdecode.scala 44:43]
  wire  _T_104 = idx_5_4; // @[dspdecode.scala 44:43]
  wire  _T_107 = idx_5_5; // @[dspdecode.scala 44:43]
  wire  busy_5 = idx_5_0 | idx_5_1 | idx_5_2 | idx_5_3 | idx_5_4 | idx_5_5; // @[dspdecode.scala 45:30]
  wire  uop_wbvld = uop_decoder_12; // @[Decodeunit.scala 13:31]
  wire [5:0] uop_wbreq = uop_decoder_37; // @[Cat.scala 30:58]
  wire  waridx_0_busyvec_0 = uop_srcreq_0_valid & io_mac_r_check_0_0_valid & uop_wbreq == io_mac_r_check_0_0_bits; // @[dspdecode.scala 44:43]
  wire  waridx_0_busyvec_1 = uop_srcreq_0_valid & io_mac_r_check_0_1_valid & uop_wbreq == io_mac_r_check_0_1_bits; // @[dspdecode.scala 44:43]
  wire  waridx_0_busyvec_2 = uop_srcreq_0_valid & io_mac_r_check_0_2_valid & uop_wbreq == io_mac_r_check_0_2_bits; // @[dspdecode.scala 44:43]
  wire  waridx_0_busyvec_3 = uop_srcreq_0_valid & io_mac_r_check_0_3_valid & uop_wbreq == io_mac_r_check_0_3_bits; // @[dspdecode.scala 44:43]
  wire  waridx_0_busyvec_4 = uop_srcreq_0_valid & io_mac_r_check_0_4_valid & uop_wbreq == io_mac_r_check_0_4_bits; // @[dspdecode.scala 44:43]
  wire  waridx_0_busyvec_5 = uop_srcreq_0_valid & io_mac_r_check_0_5_valid & uop_wbreq == io_mac_r_check_0_5_bits; // @[dspdecode.scala 44:43]
  wire  waridx_1_busyvec_0 = uop_srcreq_0_valid & io_mac_r_check_1_0_valid & uop_wbreq == io_mac_r_check_1_0_bits; // @[dspdecode.scala 44:43]
  wire  waridx_1_busyvec_1 = uop_srcreq_0_valid & io_mac_r_check_1_1_valid & uop_wbreq == io_mac_r_check_1_1_bits; // @[dspdecode.scala 44:43]
  wire  waridx_1_busyvec_2 = uop_srcreq_0_valid & io_mac_r_check_1_2_valid & uop_wbreq == io_mac_r_check_1_2_bits; // @[dspdecode.scala 44:43]
  wire  waridx_1_busyvec_3 = uop_srcreq_0_valid & io_mac_r_check_1_3_valid & uop_wbreq == io_mac_r_check_1_3_bits; // @[dspdecode.scala 44:43]
  wire  waridx_1_busyvec_4 = uop_srcreq_0_valid & io_mac_r_check_1_4_valid & uop_wbreq == io_mac_r_check_1_4_bits; // @[dspdecode.scala 44:43]
  wire  waridx_1_busyvec_5 = uop_srcreq_0_valid & io_mac_r_check_1_5_valid & uop_wbreq == io_mac_r_check_1_5_bits; // @[dspdecode.scala 44:43]
  wire  waridx_2_busyvec_0 = uop_srcreq_0_valid & io_mac_r_check_2_0_valid & uop_wbreq == io_mac_r_check_2_0_bits; // @[dspdecode.scala 44:43]
  wire  waridx_2_busyvec_1 = uop_srcreq_0_valid & io_mac_r_check_2_1_valid & uop_wbreq == io_mac_r_check_2_1_bits; // @[dspdecode.scala 44:43]
  wire  waridx_2_busyvec_2 = uop_srcreq_0_valid & io_mac_r_check_2_2_valid & uop_wbreq == io_mac_r_check_2_2_bits; // @[dspdecode.scala 44:43]
  wire  waridx_2_busyvec_3 = uop_srcreq_0_valid & io_mac_r_check_2_3_valid & uop_wbreq == io_mac_r_check_2_3_bits; // @[dspdecode.scala 44:43]
  wire  waridx_2_busyvec_4 = uop_srcreq_0_valid & io_mac_r_check_2_4_valid & uop_wbreq == io_mac_r_check_2_4_bits; // @[dspdecode.scala 44:43]
  wire  waridx_2_busyvec_5 = uop_srcreq_0_valid & io_mac_r_check_2_5_valid & uop_wbreq == io_mac_r_check_2_5_bits; // @[dspdecode.scala 44:43]
  wire  waridx_3_busyvec_0 = uop_srcreq_0_valid & io_mac_r_check_3_0_valid & uop_wbreq == io_mac_r_check_3_0_bits; // @[dspdecode.scala 44:43]
  wire  waridx_3_busyvec_1 = uop_srcreq_0_valid & io_mac_r_check_3_1_valid & uop_wbreq == io_mac_r_check_3_1_bits; // @[dspdecode.scala 44:43]
  wire  waridx_3_busyvec_2 = uop_srcreq_0_valid & io_mac_r_check_3_2_valid & uop_wbreq == io_mac_r_check_3_2_bits; // @[dspdecode.scala 44:43]
  wire  waridx_3_busyvec_3 = uop_srcreq_0_valid & io_mac_r_check_3_3_valid & uop_wbreq == io_mac_r_check_3_3_bits; // @[dspdecode.scala 44:43]
  wire  waridx_3_busyvec_4 = uop_srcreq_0_valid & io_mac_r_check_3_4_valid & uop_wbreq == io_mac_r_check_3_4_bits; // @[dspdecode.scala 44:43]
  wire  waridx_3_busyvec_5 = uop_srcreq_0_valid & io_mac_r_check_3_5_valid & uop_wbreq == io_mac_r_check_3_5_bits; // @[dspdecode.scala 44:43]
  wire  waridx_4_busyvec_0 = uop_srcreq_0_valid & io_mac_r_check_4_0_valid & uop_wbreq == io_mac_r_check_4_0_bits; // @[dspdecode.scala 44:43]
  wire  waridx_4_busyvec_1 = uop_srcreq_0_valid & io_mac_r_check_4_1_valid & uop_wbreq == io_mac_r_check_4_1_bits; // @[dspdecode.scala 44:43]
  wire  waridx_4_busyvec_2 = uop_srcreq_0_valid & io_mac_r_check_4_2_valid & uop_wbreq == io_mac_r_check_4_2_bits; // @[dspdecode.scala 44:43]
  wire  waridx_4_busyvec_3 = uop_srcreq_0_valid & io_mac_r_check_4_3_valid & uop_wbreq == io_mac_r_check_4_3_bits; // @[dspdecode.scala 44:43]
  wire  waridx_4_busyvec_4 = uop_srcreq_0_valid & io_mac_r_check_4_4_valid & uop_wbreq == io_mac_r_check_4_4_bits; // @[dspdecode.scala 44:43]
  wire  waridx_4_busyvec_5 = uop_srcreq_0_valid & io_mac_r_check_4_5_valid & uop_wbreq == io_mac_r_check_4_5_bits; // @[dspdecode.scala 44:43]
  wire  waridx_5_busyvec_0 = uop_srcreq_0_valid & io_cor_r_check_0_valid & uop_wbreq == io_cor_r_check_0_bits; // @[dspdecode.scala 44:43]
  wire  waridx_5_busyvec_1 = uop_srcreq_0_valid & io_cor_r_check_1_valid & uop_wbreq == io_cor_r_check_1_bits; // @[dspdecode.scala 44:43]
  wire  uop_ismacu = uop_decoder_0; // @[Decodeunit.scala 13:31]
  wire  macu_stall = uop_ismacu & ~(io_macuio_0_ready | io_macuio_1_ready | io_macuio_2_ready | io_macuio_3_ready |
    io_macuio_4_ready); // @[dspdecode.scala 108:31]
  wire [2:0] _req_port_T = io_macuio_3_ready ? 3'h3 : 3'h4; // @[Mux.scala 47:69]
  wire [2:0] _req_port_T_1 = io_macuio_2_ready ? 3'h2 : _req_port_T; // @[Mux.scala 47:69]
  wire [2:0] _req_port_T_2 = io_macuio_1_ready ? 3'h1 : _req_port_T_1; // @[Mux.scala 47:69]
  wire [2:0] req_port = io_macuio_0_ready ? 3'h0 : _req_port_T_2; // @[Mux.scala 47:69]
  wire  readwrite_en = io_exuempty_0 & io_exuempty_1 & io_exuempty_2 & io_exuempty_3 & io_exuempty_4 & io_exuempty_5; // @[dspdecode.scala 121:43]
  wire  uop_isread = uop_decoder_2; // @[Decodeunit.scala 12:125]
  wire [31:0] _io_writerf_bits_2_out_T_2 = io_coef_in_mainch_ch0_inputsel == 3'h1 ? io_din_bits_1 : 32'h0; // @[dspdecode.scala 129:10]
  wire [31:0] _io_writerf_bits_3_out_T_2 = io_coef_in_mainch_ch1_inputsel == 3'h1 ? io_din_bits_1 : 32'h0; // @[dspdecode.scala 129:10]
  wire  uop_iswrite = uop_decoder_3; // @[Decodeunit.scala 12:125]
  wire  uop_iscoru = uop_decoder_1; // @[Decodeunit.scala 13:31]
  wire  _stall_T_2 = uop_iscoru & ~io_coruio_ready; // @[dspdecode.scala 145:16]
  wire  _stall_T_3 = uop_ismacu & macu_stall | _stall_T_2; // @[dspdecode.scala 144:40]
  wire  _stall_T_6 = _uop_decoder_bit_T_113 & ~(readwrite_en & io_din_valid); // @[dspdecode.scala 146:16]
  wire  _stall_T_7 = _stall_T_3 | _stall_T_6; // @[dspdecode.scala 145:36]
  wire  _stall_T_10 = _uop_decoder_bit_T_115 & ~(readwrite_en & io_dout_ready); // @[dspdecode.scala 147:17]
  wire  stall = _stall_T_7 | _stall_T_10; // @[dspdecode.scala 146:51]
  wire [5:0] _instcnt_T_2 = instcnt + 6'h1; // @[dspdecode.scala 155:56]
  wire  uop_cortype = uop_decoder_4; // @[Decodeunit.scala 12:125]
  wire [2:0] uop_vlen = uop_decoder_5; // @[Cat.scala 30:58]
  wire  uop_select = uop_decoder_6; // @[Decodeunit.scala 13:31]
  wire  uop_loop = uop_decoder_7; // @[Decodeunit.scala 13:31]
  wire  uop_drc = uop_decoder_8; // @[Decodeunit.scala 13:31]
  wire  uop_pow = uop_decoder_9; // @[Decodeunit.scala 13:31]
  wire  uop_drcgain = uop_decoder_10; // @[Decodeunit.scala 13:31]
  wire  uop_drcnum = uop_decoder_11; // @[Decodeunit.scala 12:125]
  wire  uop_srcreq_0_isgroup = 1'h0; // @[dspdecode.scala 76:17 decode.scala 116:42]
  wire  _busy_T_4 = busy; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_0_busy = busy; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_0_wkupidx_0 = idx__0; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_0_wkupidx_1 = idx__1; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_0_wkupidx_2 = idx__2; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_0_wkupidx_3 = idx__3; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_0_wkupidx_4 = idx__4; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_0_wkupidx_5 = idx__5; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_1_isgroup = uop_decoder_17; // @[Decodeunit.scala 13:31]
  wire  _busy_T_9 = busy_1; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_1_busy = busy_1; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_1_wkupidx_0 = idx_1_0; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_1_wkupidx_1 = idx_1_1; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_1_wkupidx_2 = idx_1_2; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_1_wkupidx_3 = idx_1_3; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_1_wkupidx_4 = idx_1_4; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_1_wkupidx_5 = idx_1_5; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_2_isgroup = uop_decoder_21; // @[Decodeunit.scala 13:31]
  wire  _busy_T_14 = busy_2; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_2_busy = busy_2; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_2_wkupidx_0 = idx_2_0; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_2_wkupidx_1 = idx_2_1; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_2_wkupidx_2 = idx_2_2; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_2_wkupidx_3 = idx_2_3; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_2_wkupidx_4 = idx_2_4; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_2_wkupidx_5 = idx_2_5; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_3_isgroup = uop_decoder_25; // @[Decodeunit.scala 13:31]
  wire  _busy_T_19 = busy_3; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_3_busy = busy_3; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_3_wkupidx_0 = idx_3_0; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_3_wkupidx_1 = idx_3_1; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_3_wkupidx_2 = idx_3_2; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_3_wkupidx_3 = idx_3_3; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_3_wkupidx_4 = idx_3_4; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_3_wkupidx_5 = idx_3_5; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_4_isgroup = 1'h1; // @[Decodeunit.scala 13:31]
  wire  _busy_T_24 = busy_4; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_4_busy = busy_4; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_4_wkupidx_0 = idx_4_0; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_4_wkupidx_1 = idx_4_1; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_4_wkupidx_2 = idx_4_2; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_4_wkupidx_3 = idx_4_3; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_4_wkupidx_4 = idx_4_4; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_4_wkupidx_5 = idx_4_5; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_5_isgroup = uop_decoder_33; // @[Decodeunit.scala 13:31]
  wire  _busy_T_29 = busy_5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_5_busy = busy_5; // @[dspdecode.scala 45:30]
  wire  uop_srcreq_5_wkupidx_0 = idx_5_0; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_5_wkupidx_1 = idx_5_1; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_5_wkupidx_2 = idx_5_2; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_5_wkupidx_3 = idx_5_3; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_5_wkupidx_4 = idx_5_4; // @[dspdecode.scala 44:43]
  wire  uop_srcreq_5_wkupidx_5 = idx_5_5; // @[dspdecode.scala 44:43]
  assign io_din_ready = _uop_decoder_bit_T_113 & readwrite_en & io_din_valid; // @[dspdecode.scala 138:46]
  assign io_dout_valid = _uop_decoder_bit_T_115 & readwrite_en; // @[dspdecode.scala 140:32]
  assign io_dout_bits_0 = io_readrf_0; // @[dspdecode.scala 141:16]
  assign io_dout_bits_1 = io_readrf_1; // @[dspdecode.scala 141:16]
  assign io_macuio_0_valid = 3'h0 == req_port & uop_ismacu; // @[dspdecode.scala 110:29 dspdecode.scala 110:29 dspdecode.scala 101:24]
  assign io_macuio_0_bits_vlen = uop_vlen; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_select = uop_select; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_drc = uop_drc; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_pow = uop_pow; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_loop = uop_loop; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_drcgain = uop_drcgain; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_drcnum = _uop_decoder_T_21; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_valid = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_isgroup = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_idx = uop_srcreq_0_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_busy = _busy_T_4; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_wkupidx_0 = _T_2; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_wkupidx_1 = _T_5; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_wkupidx_2 = _T_8; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_wkupidx_3 = _T_11; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_wkupidx_4 = _T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_0_wkupidx_5 = _T_17; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_valid = uop_srcreq_1_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_isgroup = uop_srcreq_1_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_idx = uop_srcreq_1_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_busy = _busy_T_9; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_wkupidx_0 = _T_20; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_wkupidx_1 = _T_23; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_wkupidx_2 = _T_26; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_wkupidx_3 = _T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_wkupidx_4 = _T_32; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_1_wkupidx_5 = _T_35; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_valid = uop_srcreq_2_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_isgroup = uop_srcreq_2_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_idx = uop_srcreq_2_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_busy = _busy_T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_wkupidx_0 = _T_38; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_wkupidx_1 = _T_41; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_wkupidx_2 = _T_44; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_wkupidx_3 = _T_47; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_wkupidx_4 = _T_50; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_2_wkupidx_5 = _T_53; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_valid = uop_srcreq_3_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_isgroup = uop_srcreq_3_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_idx = uop_srcreq_3_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_busy = _busy_T_19; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_wkupidx_0 = _T_56; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_wkupidx_1 = _T_59; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_wkupidx_2 = _T_62; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_wkupidx_3 = _T_65; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_wkupidx_4 = _T_68; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_3_wkupidx_5 = _T_71; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_valid = uop_srcreq_4_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_isgroup = _uop_decoder_T_337; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_idx = uop_srcreq_4_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_busy = _busy_T_24; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_wkupidx_0 = _T_74; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_wkupidx_1 = _T_77; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_wkupidx_2 = _T_80; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_wkupidx_3 = _T_83; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_wkupidx_4 = _T_86; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_4_wkupidx_5 = _T_89; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_valid = uop_srcreq_5_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_isgroup = uop_srcreq_5_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_iscoef = uop_srcreq_5_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_idx = uop_srcreq_5_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_busy = _busy_T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_wkupidx_0 = _T_92; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_wkupidx_1 = _T_95; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_wkupidx_2 = _T_98; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_wkupidx_3 = _T_101; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_wkupidx_4 = _T_104; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_srcreq_5_wkupidx_5 = _T_107; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_wbvld = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_wbreq = uop_wbreq; // @[dspdecode.scala 102:23]
  assign io_macuio_0_bits_waridx_0 = waridx_1_busyvec_0 | waridx_1_busyvec_1 | waridx_1_busyvec_2 | waridx_1_busyvec_3
     | waridx_1_busyvec_4 | waridx_1_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_0_bits_waridx_1 = waridx_2_busyvec_0 | waridx_2_busyvec_1 | waridx_2_busyvec_2 | waridx_2_busyvec_3
     | waridx_2_busyvec_4 | waridx_2_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_0_bits_waridx_2 = waridx_3_busyvec_0 | waridx_3_busyvec_1 | waridx_3_busyvec_2 | waridx_3_busyvec_3
     | waridx_3_busyvec_4 | waridx_3_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_0_bits_waridx_3 = waridx_4_busyvec_0 | waridx_4_busyvec_1 | waridx_4_busyvec_2 | waridx_4_busyvec_3
     | waridx_4_busyvec_4 | waridx_4_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_0_bits_waridx_4 = waridx_5_busyvec_0 | waridx_5_busyvec_1; // @[dspdecode.scala 45:30]
  assign io_macuio_0_bits_wawidx_0 = uop_srcreq_0_valid & io_wd_check_1_valid & uop_wbreq == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_0_bits_wawidx_1 = uop_srcreq_0_valid & io_wd_check_2_valid & uop_wbreq == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_0_bits_wawidx_2 = uop_srcreq_0_valid & io_wd_check_3_valid & uop_wbreq == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_0_bits_wawidx_3 = uop_srcreq_0_valid & io_wd_check_4_valid & uop_wbreq == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_0_bits_wawidx_4 = uop_srcreq_0_valid & io_wd_check_5_valid & uop_wbreq == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_1_valid = 3'h1 == req_port & uop_ismacu; // @[dspdecode.scala 110:29 dspdecode.scala 110:29 dspdecode.scala 101:24]
  assign io_macuio_1_bits_vlen = uop_vlen; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_select = uop_select; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_drc = uop_drc; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_pow = uop_pow; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_loop = uop_loop; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_drcgain = uop_drcgain; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_drcnum = _uop_decoder_T_21; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_valid = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_isgroup = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_idx = uop_srcreq_0_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_busy = _busy_T_4; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_wkupidx_0 = _T_2; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_wkupidx_1 = _T_5; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_wkupidx_2 = _T_8; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_wkupidx_3 = _T_11; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_wkupidx_4 = _T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_0_wkupidx_5 = _T_17; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_valid = uop_srcreq_1_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_isgroup = uop_srcreq_1_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_idx = uop_srcreq_1_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_busy = _busy_T_9; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_wkupidx_0 = _T_20; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_wkupidx_1 = _T_23; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_wkupidx_2 = _T_26; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_wkupidx_3 = _T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_wkupidx_4 = _T_32; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_1_wkupidx_5 = _T_35; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_valid = uop_srcreq_2_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_isgroup = uop_srcreq_2_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_idx = uop_srcreq_2_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_busy = _busy_T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_wkupidx_0 = _T_38; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_wkupidx_1 = _T_41; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_wkupidx_2 = _T_44; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_wkupidx_3 = _T_47; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_wkupidx_4 = _T_50; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_2_wkupidx_5 = _T_53; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_valid = uop_srcreq_3_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_isgroup = uop_srcreq_3_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_idx = uop_srcreq_3_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_busy = _busy_T_19; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_wkupidx_0 = _T_56; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_wkupidx_1 = _T_59; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_wkupidx_2 = _T_62; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_wkupidx_3 = _T_65; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_wkupidx_4 = _T_68; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_3_wkupidx_5 = _T_71; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_valid = uop_srcreq_4_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_isgroup = _uop_decoder_T_337; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_idx = uop_srcreq_4_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_busy = _busy_T_24; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_wkupidx_0 = _T_74; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_wkupidx_1 = _T_77; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_wkupidx_2 = _T_80; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_wkupidx_3 = _T_83; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_wkupidx_4 = _T_86; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_4_wkupidx_5 = _T_89; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_valid = uop_srcreq_5_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_isgroup = uop_srcreq_5_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_iscoef = uop_srcreq_5_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_idx = uop_srcreq_5_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_busy = _busy_T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_wkupidx_0 = _T_92; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_wkupidx_1 = _T_95; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_wkupidx_2 = _T_98; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_wkupidx_3 = _T_101; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_wkupidx_4 = _T_104; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_srcreq_5_wkupidx_5 = _T_107; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_wbvld = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_wbreq = uop_wbreq; // @[dspdecode.scala 102:23]
  assign io_macuio_1_bits_waridx_0 = waridx_0_busyvec_0 | waridx_0_busyvec_1 | waridx_0_busyvec_2 | waridx_0_busyvec_3
     | waridx_0_busyvec_4 | waridx_0_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_1_bits_waridx_1 = waridx_2_busyvec_0 | waridx_2_busyvec_1 | waridx_2_busyvec_2 | waridx_2_busyvec_3
     | waridx_2_busyvec_4 | waridx_2_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_1_bits_waridx_2 = waridx_3_busyvec_0 | waridx_3_busyvec_1 | waridx_3_busyvec_2 | waridx_3_busyvec_3
     | waridx_3_busyvec_4 | waridx_3_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_1_bits_waridx_3 = waridx_4_busyvec_0 | waridx_4_busyvec_1 | waridx_4_busyvec_2 | waridx_4_busyvec_3
     | waridx_4_busyvec_4 | waridx_4_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_1_bits_waridx_4 = waridx_5_busyvec_0 | waridx_5_busyvec_1; // @[dspdecode.scala 45:30]
  assign io_macuio_1_bits_wawidx_0 = uop_srcreq_0_valid & io_wd_check_0_valid & uop_wbreq == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_1_bits_wawidx_1 = uop_srcreq_0_valid & io_wd_check_2_valid & uop_wbreq == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_1_bits_wawidx_2 = uop_srcreq_0_valid & io_wd_check_3_valid & uop_wbreq == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_1_bits_wawidx_3 = uop_srcreq_0_valid & io_wd_check_4_valid & uop_wbreq == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_1_bits_wawidx_4 = uop_srcreq_0_valid & io_wd_check_5_valid & uop_wbreq == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_2_valid = 3'h2 == req_port & uop_ismacu; // @[dspdecode.scala 110:29 dspdecode.scala 110:29 dspdecode.scala 101:24]
  assign io_macuio_2_bits_vlen = uop_vlen; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_select = uop_select; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_drc = uop_drc; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_pow = uop_pow; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_loop = uop_loop; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_drcgain = uop_drcgain; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_drcnum = _uop_decoder_T_21; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_valid = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_isgroup = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_idx = uop_srcreq_0_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_busy = _busy_T_4; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_wkupidx_0 = _T_2; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_wkupidx_1 = _T_5; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_wkupidx_2 = _T_8; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_wkupidx_3 = _T_11; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_wkupidx_4 = _T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_0_wkupidx_5 = _T_17; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_valid = uop_srcreq_1_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_isgroup = uop_srcreq_1_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_idx = uop_srcreq_1_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_busy = _busy_T_9; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_wkupidx_0 = _T_20; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_wkupidx_1 = _T_23; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_wkupidx_2 = _T_26; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_wkupidx_3 = _T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_wkupidx_4 = _T_32; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_1_wkupidx_5 = _T_35; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_valid = uop_srcreq_2_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_isgroup = uop_srcreq_2_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_idx = uop_srcreq_2_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_busy = _busy_T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_wkupidx_0 = _T_38; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_wkupidx_1 = _T_41; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_wkupidx_2 = _T_44; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_wkupidx_3 = _T_47; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_wkupidx_4 = _T_50; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_2_wkupidx_5 = _T_53; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_valid = uop_srcreq_3_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_isgroup = uop_srcreq_3_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_idx = uop_srcreq_3_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_busy = _busy_T_19; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_wkupidx_0 = _T_56; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_wkupidx_1 = _T_59; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_wkupidx_2 = _T_62; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_wkupidx_3 = _T_65; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_wkupidx_4 = _T_68; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_3_wkupidx_5 = _T_71; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_valid = uop_srcreq_4_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_isgroup = _uop_decoder_T_337; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_idx = uop_srcreq_4_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_busy = _busy_T_24; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_wkupidx_0 = _T_74; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_wkupidx_1 = _T_77; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_wkupidx_2 = _T_80; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_wkupidx_3 = _T_83; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_wkupidx_4 = _T_86; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_4_wkupidx_5 = _T_89; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_valid = uop_srcreq_5_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_isgroup = uop_srcreq_5_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_iscoef = uop_srcreq_5_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_idx = uop_srcreq_5_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_busy = _busy_T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_wkupidx_0 = _T_92; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_wkupidx_1 = _T_95; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_wkupidx_2 = _T_98; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_wkupidx_3 = _T_101; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_wkupidx_4 = _T_104; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_srcreq_5_wkupidx_5 = _T_107; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_wbvld = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_wbreq = uop_wbreq; // @[dspdecode.scala 102:23]
  assign io_macuio_2_bits_waridx_0 = waridx_0_busyvec_0 | waridx_0_busyvec_1 | waridx_0_busyvec_2 | waridx_0_busyvec_3
     | waridx_0_busyvec_4 | waridx_0_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_2_bits_waridx_1 = waridx_1_busyvec_0 | waridx_1_busyvec_1 | waridx_1_busyvec_2 | waridx_1_busyvec_3
     | waridx_1_busyvec_4 | waridx_1_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_2_bits_waridx_2 = waridx_3_busyvec_0 | waridx_3_busyvec_1 | waridx_3_busyvec_2 | waridx_3_busyvec_3
     | waridx_3_busyvec_4 | waridx_3_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_2_bits_waridx_3 = waridx_4_busyvec_0 | waridx_4_busyvec_1 | waridx_4_busyvec_2 | waridx_4_busyvec_3
     | waridx_4_busyvec_4 | waridx_4_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_2_bits_waridx_4 = waridx_5_busyvec_0 | waridx_5_busyvec_1; // @[dspdecode.scala 45:30]
  assign io_macuio_2_bits_wawidx_0 = uop_srcreq_0_valid & io_wd_check_0_valid & uop_wbreq == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_2_bits_wawidx_1 = uop_srcreq_0_valid & io_wd_check_1_valid & uop_wbreq == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_2_bits_wawidx_2 = uop_srcreq_0_valid & io_wd_check_3_valid & uop_wbreq == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_2_bits_wawidx_3 = uop_srcreq_0_valid & io_wd_check_4_valid & uop_wbreq == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_2_bits_wawidx_4 = uop_srcreq_0_valid & io_wd_check_5_valid & uop_wbreq == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_3_valid = 3'h3 == req_port & uop_ismacu; // @[dspdecode.scala 110:29 dspdecode.scala 110:29 dspdecode.scala 101:24]
  assign io_macuio_3_bits_vlen = uop_vlen; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_select = uop_select; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_drc = uop_drc; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_pow = uop_pow; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_loop = uop_loop; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_drcgain = uop_drcgain; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_drcnum = _uop_decoder_T_21; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_valid = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_isgroup = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_idx = uop_srcreq_0_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_busy = _busy_T_4; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_wkupidx_0 = _T_2; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_wkupidx_1 = _T_5; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_wkupidx_2 = _T_8; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_wkupidx_3 = _T_11; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_wkupidx_4 = _T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_0_wkupidx_5 = _T_17; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_valid = uop_srcreq_1_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_isgroup = uop_srcreq_1_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_idx = uop_srcreq_1_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_busy = _busy_T_9; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_wkupidx_0 = _T_20; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_wkupidx_1 = _T_23; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_wkupidx_2 = _T_26; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_wkupidx_3 = _T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_wkupidx_4 = _T_32; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_1_wkupidx_5 = _T_35; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_valid = uop_srcreq_2_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_isgroup = uop_srcreq_2_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_idx = uop_srcreq_2_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_busy = _busy_T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_wkupidx_0 = _T_38; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_wkupidx_1 = _T_41; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_wkupidx_2 = _T_44; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_wkupidx_3 = _T_47; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_wkupidx_4 = _T_50; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_2_wkupidx_5 = _T_53; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_valid = uop_srcreq_3_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_isgroup = uop_srcreq_3_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_idx = uop_srcreq_3_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_busy = _busy_T_19; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_wkupidx_0 = _T_56; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_wkupidx_1 = _T_59; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_wkupidx_2 = _T_62; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_wkupidx_3 = _T_65; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_wkupidx_4 = _T_68; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_3_wkupidx_5 = _T_71; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_valid = uop_srcreq_4_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_isgroup = _uop_decoder_T_337; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_idx = uop_srcreq_4_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_busy = _busy_T_24; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_wkupidx_0 = _T_74; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_wkupidx_1 = _T_77; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_wkupidx_2 = _T_80; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_wkupidx_3 = _T_83; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_wkupidx_4 = _T_86; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_4_wkupidx_5 = _T_89; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_valid = uop_srcreq_5_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_isgroup = uop_srcreq_5_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_iscoef = uop_srcreq_5_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_idx = uop_srcreq_5_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_busy = _busy_T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_wkupidx_0 = _T_92; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_wkupidx_1 = _T_95; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_wkupidx_2 = _T_98; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_wkupidx_3 = _T_101; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_wkupidx_4 = _T_104; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_srcreq_5_wkupidx_5 = _T_107; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_wbvld = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_wbreq = uop_wbreq; // @[dspdecode.scala 102:23]
  assign io_macuio_3_bits_waridx_0 = waridx_0_busyvec_0 | waridx_0_busyvec_1 | waridx_0_busyvec_2 | waridx_0_busyvec_3
     | waridx_0_busyvec_4 | waridx_0_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_3_bits_waridx_1 = waridx_1_busyvec_0 | waridx_1_busyvec_1 | waridx_1_busyvec_2 | waridx_1_busyvec_3
     | waridx_1_busyvec_4 | waridx_1_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_3_bits_waridx_2 = waridx_2_busyvec_0 | waridx_2_busyvec_1 | waridx_2_busyvec_2 | waridx_2_busyvec_3
     | waridx_2_busyvec_4 | waridx_2_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_3_bits_waridx_3 = waridx_4_busyvec_0 | waridx_4_busyvec_1 | waridx_4_busyvec_2 | waridx_4_busyvec_3
     | waridx_4_busyvec_4 | waridx_4_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_3_bits_waridx_4 = waridx_5_busyvec_0 | waridx_5_busyvec_1; // @[dspdecode.scala 45:30]
  assign io_macuio_3_bits_wawidx_0 = uop_srcreq_0_valid & io_wd_check_0_valid & uop_wbreq == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_3_bits_wawidx_1 = uop_srcreq_0_valid & io_wd_check_1_valid & uop_wbreq == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_3_bits_wawidx_2 = uop_srcreq_0_valid & io_wd_check_2_valid & uop_wbreq == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_3_bits_wawidx_3 = uop_srcreq_0_valid & io_wd_check_4_valid & uop_wbreq == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_3_bits_wawidx_4 = uop_srcreq_0_valid & io_wd_check_5_valid & uop_wbreq == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_4_valid = 3'h4 == req_port & uop_ismacu; // @[dspdecode.scala 110:29 dspdecode.scala 110:29 dspdecode.scala 101:24]
  assign io_macuio_4_bits_vlen = uop_vlen; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_select = uop_select; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_drc = uop_drc; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_pow = uop_pow; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_loop = uop_loop; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_drcgain = uop_drcgain; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_drcnum = _uop_decoder_T_21; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_valid = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_isgroup = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_idx = uop_srcreq_0_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_busy = _busy_T_4; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_wkupidx_0 = _T_2; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_wkupidx_1 = _T_5; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_wkupidx_2 = _T_8; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_wkupidx_3 = _T_11; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_wkupidx_4 = _T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_0_wkupidx_5 = _T_17; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_valid = uop_srcreq_1_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_isgroup = uop_srcreq_1_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_idx = uop_srcreq_1_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_busy = _busy_T_9; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_wkupidx_0 = _T_20; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_wkupidx_1 = _T_23; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_wkupidx_2 = _T_26; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_wkupidx_3 = _T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_wkupidx_4 = _T_32; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_1_wkupidx_5 = _T_35; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_valid = uop_srcreq_2_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_isgroup = uop_srcreq_2_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_idx = uop_srcreq_2_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_busy = _busy_T_14; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_wkupidx_0 = _T_38; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_wkupidx_1 = _T_41; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_wkupidx_2 = _T_44; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_wkupidx_3 = _T_47; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_wkupidx_4 = _T_50; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_2_wkupidx_5 = _T_53; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_valid = uop_srcreq_3_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_isgroup = uop_srcreq_3_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_idx = uop_srcreq_3_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_busy = _busy_T_19; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_wkupidx_0 = _T_56; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_wkupidx_1 = _T_59; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_wkupidx_2 = _T_62; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_wkupidx_3 = _T_65; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_wkupidx_4 = _T_68; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_3_wkupidx_5 = _T_71; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_valid = uop_srcreq_4_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_isgroup = _uop_decoder_T_337; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_iscoef = uop_srcreq_0_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_idx = uop_srcreq_4_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_busy = _busy_T_24; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_wkupidx_0 = _T_74; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_wkupidx_1 = _T_77; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_wkupidx_2 = _T_80; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_wkupidx_3 = _T_83; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_wkupidx_4 = _T_86; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_4_wkupidx_5 = _T_89; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_valid = uop_srcreq_5_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_isgroup = uop_srcreq_5_isgroup; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_iscoef = uop_srcreq_5_iscoef; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_idx = uop_srcreq_5_idx; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_busy = _busy_T_29; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_wkupidx_0 = _T_92; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_wkupidx_1 = _T_95; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_wkupidx_2 = _T_98; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_wkupidx_3 = _T_101; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_wkupidx_4 = _T_104; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_srcreq_5_wkupidx_5 = _T_107; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_wbvld = uop_srcreq_0_valid; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_wbreq = uop_wbreq; // @[dspdecode.scala 102:23]
  assign io_macuio_4_bits_waridx_0 = waridx_0_busyvec_0 | waridx_0_busyvec_1 | waridx_0_busyvec_2 | waridx_0_busyvec_3
     | waridx_0_busyvec_4 | waridx_0_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_4_bits_waridx_1 = waridx_1_busyvec_0 | waridx_1_busyvec_1 | waridx_1_busyvec_2 | waridx_1_busyvec_3
     | waridx_1_busyvec_4 | waridx_1_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_4_bits_waridx_2 = waridx_2_busyvec_0 | waridx_2_busyvec_1 | waridx_2_busyvec_2 | waridx_2_busyvec_3
     | waridx_2_busyvec_4 | waridx_2_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_4_bits_waridx_3 = waridx_3_busyvec_0 | waridx_3_busyvec_1 | waridx_3_busyvec_2 | waridx_3_busyvec_3
     | waridx_3_busyvec_4 | waridx_3_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_macuio_4_bits_waridx_4 = waridx_5_busyvec_0 | waridx_5_busyvec_1; // @[dspdecode.scala 45:30]
  assign io_macuio_4_bits_wawidx_0 = uop_srcreq_0_valid & io_wd_check_0_valid & uop_wbreq == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_4_bits_wawidx_1 = uop_srcreq_0_valid & io_wd_check_1_valid & uop_wbreq == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_4_bits_wawidx_2 = uop_srcreq_0_valid & io_wd_check_2_valid & uop_wbreq == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_4_bits_wawidx_3 = uop_srcreq_0_valid & io_wd_check_3_valid & uop_wbreq == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  assign io_macuio_4_bits_wawidx_4 = uop_srcreq_0_valid & io_wd_check_5_valid & uop_wbreq == io_wd_check_5_bits; // @[dspdecode.scala 44:43]
  assign io_coruio_valid = uop_iscoru; // @[dspdecode.scala 118:19]
  assign io_coruio_bits_cortype = _uop_decoder_T_1; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_valid = uop_srcreq_0_valid; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_idx = uop_srcreq_0_idx; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_busy = _busy_T_4; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_wkupidx_0 = _T_2; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_wkupidx_1 = _T_5; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_wkupidx_2 = _T_8; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_wkupidx_3 = _T_11; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_wkupidx_4 = _T_14; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_0_wkupidx_5 = _T_17; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_valid = uop_srcreq_5_valid; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_idx = uop_srcreq_5_idx; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_busy = _busy_T_29; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_wkupidx_0 = _T_92; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_wkupidx_1 = _T_95; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_wkupidx_2 = _T_98; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_wkupidx_3 = _T_101; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_wkupidx_4 = _T_104; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_srcreq_1_wkupidx_5 = _T_107; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_wbvld = uop_srcreq_0_valid; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_wbreq = uop_wbreq; // @[dspdecode.scala 115:18]
  assign io_coruio_bits_waridx_0 = waridx_0_busyvec_0 | waridx_0_busyvec_1 | waridx_0_busyvec_2 | waridx_0_busyvec_3 |
    waridx_0_busyvec_4 | waridx_0_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_coruio_bits_waridx_1 = waridx_1_busyvec_0 | waridx_1_busyvec_1 | waridx_1_busyvec_2 | waridx_1_busyvec_3 |
    waridx_1_busyvec_4 | waridx_1_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_coruio_bits_waridx_2 = waridx_2_busyvec_0 | waridx_2_busyvec_1 | waridx_2_busyvec_2 | waridx_2_busyvec_3 |
    waridx_2_busyvec_4 | waridx_2_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_coruio_bits_waridx_3 = waridx_3_busyvec_0 | waridx_3_busyvec_1 | waridx_3_busyvec_2 | waridx_3_busyvec_3 |
    waridx_3_busyvec_4 | waridx_3_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_coruio_bits_waridx_4 = waridx_4_busyvec_0 | waridx_4_busyvec_1 | waridx_4_busyvec_2 | waridx_4_busyvec_3 |
    waridx_4_busyvec_4 | waridx_4_busyvec_5; // @[dspdecode.scala 45:30]
  assign io_coruio_bits_wawidx_0 = uop_srcreq_0_valid & io_wd_check_0_valid & uop_wbreq == io_wd_check_0_bits; // @[dspdecode.scala 44:43]
  assign io_coruio_bits_wawidx_1 = uop_srcreq_0_valid & io_wd_check_1_valid & uop_wbreq == io_wd_check_1_bits; // @[dspdecode.scala 44:43]
  assign io_coruio_bits_wawidx_2 = uop_srcreq_0_valid & io_wd_check_2_valid & uop_wbreq == io_wd_check_2_bits; // @[dspdecode.scala 44:43]
  assign io_coruio_bits_wawidx_3 = uop_srcreq_0_valid & io_wd_check_3_valid & uop_wbreq == io_wd_check_3_bits; // @[dspdecode.scala 44:43]
  assign io_coruio_bits_wawidx_4 = uop_srcreq_0_valid & io_wd_check_4_valid & uop_wbreq == io_wd_check_4_bits; // @[dspdecode.scala 44:43]
  assign io_writerf_valid = readwrite_en & _uop_decoder_bit_T_113 & io_din_valid; // @[dspdecode.scala 133:50]
  assign io_writerf_bits_0 = io_din_bits_0; // @[dspdecode.scala 134:22]
  assign io_writerf_bits_1 = io_din_bits_1; // @[dspdecode.scala 135:22]
  assign io_writerf_bits_2 = io_coef_in_mainch_ch0_inputsel == 3'h0 ? io_din_bits_0 : _io_writerf_bits_2_out_T_2; // @[dspdecode.scala 128:15]
  assign io_writerf_bits_3 = io_coef_in_mainch_ch1_inputsel == 3'h0 ? io_din_bits_0 : _io_writerf_bits_3_out_T_2; // @[dspdecode.scala 128:15]
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      instcnt <= 6'h0;
    end else if (!(stall)) begin
      if (instcnt == 6'h36) begin
        instcnt <= 6'h0;
      end else begin
        instcnt <= _instcnt_T_2;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  instcnt = _RAND_0[5:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    instcnt = 6'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile(
  input         clock,
  input         reset,
  input         io_exe_rd_0_req_isgroup,
  input         io_exe_rd_0_req_iscoef,
  input  [5:0]  io_exe_rd_0_req_idx,
  input  [2:0]  io_exe_rd_0_req_gidx,
  output [31:0] io_exe_rd_0_resp,
  input         io_exe_rd_1_req_isgroup,
  input         io_exe_rd_1_req_iscoef,
  input  [5:0]  io_exe_rd_1_req_idx,
  input  [2:0]  io_exe_rd_1_req_gidx,
  input         io_exe_rd_1_req_sel,
  output [31:0] io_exe_rd_1_resp,
  input         io_exe_rd_2_req_isgroup,
  input         io_exe_rd_2_req_iscoef,
  input  [5:0]  io_exe_rd_2_req_idx,
  input  [2:0]  io_exe_rd_2_req_gidx,
  output [31:0] io_exe_rd_2_resp,
  input         io_exe_rd_3_req_isgroup,
  input         io_exe_rd_3_req_iscoef,
  input  [5:0]  io_exe_rd_3_req_idx,
  input  [2:0]  io_exe_rd_3_req_gidx,
  input         io_exe_rd_3_req_sel,
  output [31:0] io_exe_rd_3_resp,
  input         io_exe_rd_4_req_isgroup,
  input         io_exe_rd_4_req_iscoef,
  input  [5:0]  io_exe_rd_4_req_idx,
  input  [2:0]  io_exe_rd_4_req_gidx,
  output [31:0] io_exe_rd_4_resp,
  input         io_exe_rd_5_req_isgroup,
  input         io_exe_rd_5_req_iscoef,
  input  [5:0]  io_exe_rd_5_req_idx,
  input  [2:0]  io_exe_rd_5_req_gidx,
  input         io_exe_rd_5_req_sel,
  output [31:0] io_exe_rd_5_resp,
  input         io_exe_rd_6_req_isgroup,
  input         io_exe_rd_6_req_iscoef,
  input  [5:0]  io_exe_rd_6_req_idx,
  input  [2:0]  io_exe_rd_6_req_gidx,
  output [31:0] io_exe_rd_6_resp,
  input         io_exe_rd_7_req_isgroup,
  input         io_exe_rd_7_req_iscoef,
  input  [5:0]  io_exe_rd_7_req_idx,
  input  [2:0]  io_exe_rd_7_req_gidx,
  input         io_exe_rd_7_req_sel,
  output [31:0] io_exe_rd_7_resp,
  input         io_exe_rd_8_req_isgroup,
  input         io_exe_rd_8_req_iscoef,
  input  [5:0]  io_exe_rd_8_req_idx,
  input  [2:0]  io_exe_rd_8_req_gidx,
  output [31:0] io_exe_rd_8_resp,
  input         io_exe_rd_9_req_isgroup,
  input         io_exe_rd_9_req_iscoef,
  input  [5:0]  io_exe_rd_9_req_idx,
  input  [2:0]  io_exe_rd_9_req_gidx,
  input         io_exe_rd_9_req_sel,
  output [31:0] io_exe_rd_9_resp,
  input  [5:0]  io_exe_rd_10_req_idx,
  output [31:0] io_exe_rd_10_resp,
  input  [5:0]  io_exe_rd_11_req_idx,
  output [31:0] io_exe_rd_11_resp,
  input  [31:0] io_exe_wb_0_wdata1,
  input  [31:0] io_exe_wb_0_wdata2,
  input         io_exe_wb_0_vld,
  input  [5:0]  io_exe_wb_0_gregidx,
  input  [31:0] io_exe_wb_1_wdata1,
  input  [31:0] io_exe_wb_1_wdata2,
  input         io_exe_wb_1_vld,
  input  [5:0]  io_exe_wb_1_gregidx,
  input  [31:0] io_exe_wb_2_wdata1,
  input  [31:0] io_exe_wb_2_wdata2,
  input         io_exe_wb_2_vld,
  input  [5:0]  io_exe_wb_2_gregidx,
  input  [31:0] io_exe_wb_3_wdata1,
  input  [31:0] io_exe_wb_3_wdata2,
  input         io_exe_wb_3_vld,
  input  [5:0]  io_exe_wb_3_gregidx,
  input  [31:0] io_exe_wb_4_wdata1,
  input  [31:0] io_exe_wb_4_wdata2,
  input         io_exe_wb_4_vld,
  input  [5:0]  io_exe_wb_4_gregidx,
  input  [31:0] io_exe_wb_5_wdata2,
  input         io_exe_wb_5_vld,
  input  [5:0]  io_exe_wb_5_gregidx,
  input         io_dec_wb_valid,
  input  [31:0] io_dec_wb_bits_0,
  input  [31:0] io_dec_wb_bits_1,
  input  [31:0] io_dec_wb_bits_2,
  input  [31:0] io_dec_wb_bits_3,
  output [31:0] io_dec_rd_0,
  output [31:0] io_dec_rd_1,
  input  [31:0] io_coef_in_subch_ch2mix_0,
  input  [31:0] io_coef_in_subch_ch2mix_1,
  input  [31:0] io_coef_in_subch_ch2mix_2,
  input  [31:0] io_coef_in_subch_ch2bq_0_0,
  input  [31:0] io_coef_in_subch_ch2bq_0_1,
  input  [31:0] io_coef_in_subch_ch2bq_0_2,
  input  [31:0] io_coef_in_subch_ch2bq_0_3,
  input  [31:0] io_coef_in_subch_ch2bq_0_4,
  input  [31:0] io_coef_in_subch_ch2vol,
  input         io_coef_in_subch_ch2volsel,
  input         io_coef_in_subch_ch3sel,
  input  [31:0] io_coef_in_subch_ch3mix_0,
  input  [31:0] io_coef_in_subch_ch3mix_1,
  input  [31:0] io_coef_in_subch_ch3bq_0_0,
  input  [31:0] io_coef_in_subch_ch3bq_0_1,
  input  [31:0] io_coef_in_subch_ch3bq_0_2,
  input  [31:0] io_coef_in_subch_ch3bq_0_3,
  input  [31:0] io_coef_in_subch_ch3bq_0_4,
  input  [31:0] io_coef_in_subch_ch3bq_1_0,
  input  [31:0] io_coef_in_subch_ch3bq_1_1,
  input  [31:0] io_coef_in_subch_ch3bq_1_2,
  input  [31:0] io_coef_in_subch_ch3bq_1_3,
  input  [31:0] io_coef_in_subch_ch3bq_1_4,
  input  [31:0] io_coef_in_subch_ch3vol,
  input         io_coef_in_subch_ch3volsel,
  input  [31:0] io_coef_in_subch_drc_pow_0,
  input  [31:0] io_coef_in_subch_drc_pow_1,
  input  [31:0] io_coef_in_subch_drc_smooth_0,
  input  [31:0] io_coef_in_subch_drc_smooth_1,
  input  [31:0] io_coef_in_subch_drc_smooth_2,
  input  [31:0] io_coef_in_subch_drc_smooth_3,
  input  [31:0] io_coef_in_subch_drc_ratio,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_0_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_0_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_0_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_0_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_0_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_1_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_1_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_1_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_1_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_1_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_2_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_2_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_2_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_2_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_2_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_3_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_3_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_3_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_3_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_3_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_4_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_4_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_4_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_4_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_4_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_5_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_5_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_5_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_5_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_5_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_6_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_6_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_6_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_6_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_6_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_7_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_7_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_7_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_7_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_7_4,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_8_0,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_8_1,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_8_2,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_8_3,
  input  [31:0] io_coef_in_mainch_ch0_bqcoef_8_4,
  input  [31:0] io_coef_in_mainch_ch0_inputmix_0_0,
  input  [31:0] io_coef_in_mainch_ch0_inputmix_0_1,
  input  [31:0] io_coef_in_mainch_ch0_inputmix_1_0,
  input  [31:0] io_coef_in_mainch_ch0_inputmix_1_1,
  input  [31:0] io_coef_in_mainch_ch0_vol,
  input  [31:0] io_coef_in_mainch_ch0_outputmix_0,
  input  [31:0] io_coef_in_mainch_ch0_outputmix_1,
  input  [31:0] io_coef_in_mainch_ch0_outputmix_2,
  input  [31:0] io_coef_in_mainch_ch0_prescale,
  input  [31:0] io_coef_in_mainch_ch0_postscale,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_0_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_0_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_0_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_0_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_0_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_1_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_1_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_1_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_1_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_1_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_2_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_2_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_2_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_2_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_2_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_3_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_3_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_3_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_3_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_3_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_4_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_4_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_4_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_4_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_4_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_5_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_5_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_5_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_5_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_5_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_6_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_6_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_6_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_6_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_6_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_7_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_7_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_7_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_7_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_7_4,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_8_0,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_8_1,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_8_2,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_8_3,
  input  [31:0] io_coef_in_mainch_ch1_bqcoef_8_4,
  input  [31:0] io_coef_in_mainch_ch1_inputmix_0_0,
  input  [31:0] io_coef_in_mainch_ch1_inputmix_0_1,
  input  [31:0] io_coef_in_mainch_ch1_inputmix_1_0,
  input  [31:0] io_coef_in_mainch_ch1_inputmix_1_1,
  input  [31:0] io_coef_in_mainch_ch1_vol,
  input  [31:0] io_coef_in_mainch_ch1_outputmix_0,
  input  [31:0] io_coef_in_mainch_ch1_outputmix_1,
  input  [31:0] io_coef_in_mainch_ch1_outputmix_2,
  input  [31:0] io_coef_in_mainch_drc_pow_0,
  input  [31:0] io_coef_in_mainch_drc_pow_1,
  input  [31:0] io_coef_in_mainch_drc_smooth_0,
  input  [31:0] io_coef_in_mainch_drc_smooth_1,
  input  [31:0] io_coef_in_mainch_drc_smooth_2,
  input  [31:0] io_coef_in_mainch_drc_smooth_3,
  input  [31:0] io_coef_in_mainch_drc_ratio
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_type1_data_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_0 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h0 ? io_exe_wb_0_wdata2 : reg_type1_data_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_1 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h0 ? io_exe_wb_1_wdata2 : _GEN_0; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_2 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h0 ? io_exe_wb_2_wdata2 : _GEN_1; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_3 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h0 ? io_exe_wb_3_wdata2 : _GEN_2; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_4 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h0 ? io_exe_wb_4_wdata2 : _GEN_3; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type1_data_nxt_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h0 ? io_exe_wb_5_wdata2 : _GEN_4; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type1_data_1_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_6 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1 ? io_exe_wb_0_wdata2 : reg_type1_data_1_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_7 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1 ? io_exe_wb_1_wdata2 : _GEN_6; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_8 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1 ? io_exe_wb_2_wdata2 : _GEN_7; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_9 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1 ? io_exe_wb_3_wdata2 : _GEN_8; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_10 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1 ? io_exe_wb_4_wdata2 : _GEN_9; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type1_data_nxt_1_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1 ? io_exe_wb_5_wdata2 : _GEN_10; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type1_data_2_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_12 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h2 ? io_exe_wb_0_wdata2 : reg_type1_data_2_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_13 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h2 ? io_exe_wb_1_wdata2 : _GEN_12; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_14 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h2 ? io_exe_wb_2_wdata2 : _GEN_13; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_15 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h2 ? io_exe_wb_3_wdata2 : _GEN_14; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_16 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h2 ? io_exe_wb_4_wdata2 : _GEN_15; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type1_data_nxt_2_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h2 ? io_exe_wb_5_wdata2 : _GEN_16; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type1_data_3_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_18 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h3 ? io_exe_wb_0_wdata2 : reg_type1_data_3_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_19 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h3 ? io_exe_wb_1_wdata2 : _GEN_18; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_20 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h3 ? io_exe_wb_2_wdata2 : _GEN_19; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_21 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h3 ? io_exe_wb_3_wdata2 : _GEN_20; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_22 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h3 ? io_exe_wb_4_wdata2 : _GEN_21; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type1_data_nxt_3_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h3 ? io_exe_wb_5_wdata2 : _GEN_22; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type2_data_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_28 = io_dec_wb_valid ? io_dec_wb_bits_0 : reg_type2_data_0; // @[regfile.scala 44:26 regfile.scala 45:25 regfile.scala 40:18]
  wire [31:0] _GEN_29 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h4 ? io_exe_wb_0_wdata2 : _GEN_28; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_30 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h4 ? io_exe_wb_1_wdata2 : _GEN_29; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_31 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h4 ? io_exe_wb_2_wdata2 : _GEN_30; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_32 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h4 ? io_exe_wb_3_wdata2 : _GEN_31; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_33 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h4 ? io_exe_wb_4_wdata2 : _GEN_32; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type2_data_nxt_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h4 ? io_exe_wb_5_wdata2 : _GEN_33; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type2_data_1_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_39 = io_dec_wb_valid ? io_dec_wb_bits_1 : reg_type2_data_1_0; // @[regfile.scala 44:26 regfile.scala 45:25 regfile.scala 40:18]
  wire [31:0] _GEN_40 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h5 ? io_exe_wb_0_wdata2 : _GEN_39; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_41 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h5 ? io_exe_wb_1_wdata2 : _GEN_40; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_42 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h5 ? io_exe_wb_2_wdata2 : _GEN_41; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_43 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h5 ? io_exe_wb_3_wdata2 : _GEN_42; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_44 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h5 ? io_exe_wb_4_wdata2 : _GEN_43; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type2_data_nxt_1_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h5 ? io_exe_wb_5_wdata2 : _GEN_44; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type2_data_2_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_50 = io_dec_wb_valid ? io_dec_wb_bits_2 : reg_type2_data_2_0; // @[regfile.scala 44:26 regfile.scala 45:25 regfile.scala 40:18]
  wire [31:0] _GEN_51 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h6 ? io_exe_wb_0_wdata2 : _GEN_50; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_52 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h6 ? io_exe_wb_1_wdata2 : _GEN_51; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_53 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h6 ? io_exe_wb_2_wdata2 : _GEN_52; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_54 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h6 ? io_exe_wb_3_wdata2 : _GEN_53; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_55 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h6 ? io_exe_wb_4_wdata2 : _GEN_54; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type2_data_nxt_2_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h6 ? io_exe_wb_5_wdata2 : _GEN_55; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type2_data_3_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_61 = io_dec_wb_valid ? io_dec_wb_bits_3 : reg_type2_data_3_0; // @[regfile.scala 44:26 regfile.scala 45:25 regfile.scala 40:18]
  wire [31:0] _GEN_62 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h7 ? io_exe_wb_0_wdata2 : _GEN_61; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_63 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h7 ? io_exe_wb_1_wdata2 : _GEN_62; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_64 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h7 ? io_exe_wb_2_wdata2 : _GEN_63; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_65 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h7 ? io_exe_wb_3_wdata2 : _GEN_64; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_66 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h7 ? io_exe_wb_4_wdata2 : _GEN_65; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type2_data_nxt_3_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h7 ? io_exe_wb_5_wdata2 : _GEN_66; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type3_data_0; // @[regfile.scala 21:31]
  wire [31:0] _GEN_68 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h8 ? io_exe_wb_0_wdata2 : reg_type3_data_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_69 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h8 ? io_exe_wb_1_wdata2 : _GEN_68; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_70 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h8 ? io_exe_wb_2_wdata2 : _GEN_69; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_71 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h8 ? io_exe_wb_3_wdata2 : _GEN_70; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_72 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h8 ? io_exe_wb_4_wdata2 : _GEN_71; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type3_data_nxt_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h8 ? io_exe_wb_5_wdata2 : _GEN_72; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type3_data_1_0; // @[regfile.scala 21:31]
  wire [31:0] _GEN_74 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h9 ? io_exe_wb_0_wdata2 : reg_type3_data_1_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_75 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h9 ? io_exe_wb_1_wdata2 : _GEN_74; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_76 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h9 ? io_exe_wb_2_wdata2 : _GEN_75; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_77 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h9 ? io_exe_wb_3_wdata2 : _GEN_76; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_78 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h9 ? io_exe_wb_4_wdata2 : _GEN_77; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type3_data_nxt_1_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h9 ? io_exe_wb_5_wdata2 : _GEN_78; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type4_data_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_80 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'ha ? io_exe_wb_0_wdata2 : reg_type4_data_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_81 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'ha ? io_exe_wb_1_wdata2 : _GEN_80; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_82 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'ha ? io_exe_wb_2_wdata2 : _GEN_81; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_83 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'ha ? io_exe_wb_3_wdata2 : _GEN_82; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_84 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'ha ? io_exe_wb_4_wdata2 : _GEN_83; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type4_data_nxt_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'ha ? io_exe_wb_5_wdata2 : _GEN_84; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type4_data_1_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_86 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hb ? io_exe_wb_0_wdata2 : reg_type4_data_1_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_87 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hb ? io_exe_wb_1_wdata2 : _GEN_86; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_88 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hb ? io_exe_wb_2_wdata2 : _GEN_87; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_89 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hb ? io_exe_wb_3_wdata2 : _GEN_88; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_90 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hb ? io_exe_wb_4_wdata2 : _GEN_89; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type4_data_nxt_1_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hb ? io_exe_wb_5_wdata2 : _GEN_90; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type4_data_2_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_92 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hc ? io_exe_wb_0_wdata2 : reg_type4_data_2_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_93 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hc ? io_exe_wb_1_wdata2 : _GEN_92; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_94 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hc ? io_exe_wb_2_wdata2 : _GEN_93; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_95 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hc ? io_exe_wb_3_wdata2 : _GEN_94; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_96 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hc ? io_exe_wb_4_wdata2 : _GEN_95; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type4_data_nxt_2_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hc ? io_exe_wb_5_wdata2 : _GEN_96; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type4_data_3_0; // @[regfile.scala 22:22]
  wire [31:0] _GEN_98 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hd ? io_exe_wb_0_wdata2 : reg_type4_data_3_0; // @[regfile.scala 51:64 regfile.scala 58:27 regfile.scala 40:18]
  wire [31:0] _GEN_99 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hd ? io_exe_wb_1_wdata2 : _GEN_98; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_100 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hd ? io_exe_wb_2_wdata2 : _GEN_99; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_101 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hd ? io_exe_wb_3_wdata2 : _GEN_100; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] _GEN_102 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hd ? io_exe_wb_4_wdata2 : _GEN_101; // @[regfile.scala 51:64 regfile.scala 58:27]
  wire [31:0] reg_type4_data_nxt_3_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hd ? io_exe_wb_5_wdata2 : _GEN_102; // @[regfile.scala 51:64 regfile.scala 58:27]
  reg [31:0] reg_type5_data__0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data__1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data__2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data__3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_104 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'he ? io_exe_wb_0_wdata1 : reg_type5_data__0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_105 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'he ? reg_type5_data__0 : reg_type5_data__1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_106 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'he ? io_exe_wb_0_wdata2 : reg_type5_data__2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_107 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'he ? reg_type5_data__2 : reg_type5_data__3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_108 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'he ? io_exe_wb_1_wdata1 : _GEN_104; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_109 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'he ? reg_type5_data__0 : _GEN_105; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_110 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'he ? io_exe_wb_1_wdata2 : _GEN_106; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_111 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'he ? reg_type5_data__2 : _GEN_107; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_112 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he ? io_exe_wb_2_wdata1 : _GEN_108; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_113 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he ? reg_type5_data__0 : _GEN_109; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_114 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he ? io_exe_wb_2_wdata2 : _GEN_110; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_115 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he ? reg_type5_data__2 : _GEN_111; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_116 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he ? io_exe_wb_3_wdata1 : _GEN_112; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_117 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he ? reg_type5_data__0 : _GEN_113; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_118 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he ? io_exe_wb_3_wdata2 : _GEN_114; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_119 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he ? reg_type5_data__2 : _GEN_115; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_120 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he ? io_exe_wb_4_wdata1 : _GEN_116; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_121 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he ? reg_type5_data__0 : _GEN_117; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_122 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he ? io_exe_wb_4_wdata2 : _GEN_118; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_123 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he ? reg_type5_data__2 : _GEN_119; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt__0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he ? 32'h0 : _GEN_120; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt__1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he ? reg_type5_data__0 : _GEN_121; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt__2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he ? io_exe_wb_5_wdata2 : _GEN_122; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt__3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he ? reg_type5_data__2 : _GEN_123; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_1_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_1_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_1_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_1_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_128 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hf ? io_exe_wb_0_wdata1 : reg_type5_data_1_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_129 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hf ? reg_type5_data_1_0 : reg_type5_data_1_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_130 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hf ? io_exe_wb_0_wdata2 : reg_type5_data_1_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_131 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'hf ? reg_type5_data_1_2 : reg_type5_data_1_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_132 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hf ? io_exe_wb_1_wdata1 : _GEN_128; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_133 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hf ? reg_type5_data_1_0 : _GEN_129; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_134 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hf ? io_exe_wb_1_wdata2 : _GEN_130; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_135 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'hf ? reg_type5_data_1_2 : _GEN_131; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_136 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf ? io_exe_wb_2_wdata1 : _GEN_132; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_137 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf ? reg_type5_data_1_0 : _GEN_133; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_138 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf ? io_exe_wb_2_wdata2 : _GEN_134; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_139 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf ? reg_type5_data_1_2 : _GEN_135; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_140 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf ? io_exe_wb_3_wdata1 : _GEN_136; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_141 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf ? reg_type5_data_1_0 : _GEN_137; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_142 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf ? io_exe_wb_3_wdata2 : _GEN_138; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_143 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf ? reg_type5_data_1_2 : _GEN_139; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_144 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf ? io_exe_wb_4_wdata1 : _GEN_140; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_145 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf ? reg_type5_data_1_0 : _GEN_141; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_146 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf ? io_exe_wb_4_wdata2 : _GEN_142; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_147 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf ? reg_type5_data_1_2 : _GEN_143; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_1_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf ? 32'h0 : _GEN_144; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_1_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf ? reg_type5_data_1_0 : _GEN_145; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_1_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf ? io_exe_wb_5_wdata2 : _GEN_146; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_1_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf ? reg_type5_data_1_2 : _GEN_147; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_2_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_2_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_2_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_2_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_152 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h10 ? io_exe_wb_0_wdata1 : reg_type5_data_2_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_153 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h10 ? reg_type5_data_2_0 : reg_type5_data_2_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_154 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h10 ? io_exe_wb_0_wdata2 : reg_type5_data_2_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_155 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h10 ? reg_type5_data_2_2 : reg_type5_data_2_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_156 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h10 ? io_exe_wb_1_wdata1 : _GEN_152; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_157 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h10 ? reg_type5_data_2_0 : _GEN_153; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_158 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h10 ? io_exe_wb_1_wdata2 : _GEN_154; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_159 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h10 ? reg_type5_data_2_2 : _GEN_155; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_160 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10 ? io_exe_wb_2_wdata1 : _GEN_156; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_161 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10 ? reg_type5_data_2_0 : _GEN_157; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_162 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10 ? io_exe_wb_2_wdata2 : _GEN_158; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_163 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10 ? reg_type5_data_2_2 : _GEN_159; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_164 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10 ? io_exe_wb_3_wdata1 : _GEN_160; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_165 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10 ? reg_type5_data_2_0 : _GEN_161; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_166 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10 ? io_exe_wb_3_wdata2 : _GEN_162; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_167 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10 ? reg_type5_data_2_2 : _GEN_163; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_168 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10 ? io_exe_wb_4_wdata1 : _GEN_164; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_169 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10 ? reg_type5_data_2_0 : _GEN_165; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_170 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10 ? io_exe_wb_4_wdata2 : _GEN_166; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_171 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10 ? reg_type5_data_2_2 : _GEN_167; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_2_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10 ? 32'h0 : _GEN_168; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_2_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10 ? reg_type5_data_2_0 : _GEN_169; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_2_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10 ? io_exe_wb_5_wdata2 : _GEN_170; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_2_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10 ? reg_type5_data_2_2 : _GEN_171; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_3_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_3_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_3_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_3_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_176 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h11 ? io_exe_wb_0_wdata1 : reg_type5_data_3_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_177 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h11 ? reg_type5_data_3_0 : reg_type5_data_3_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_178 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h11 ? io_exe_wb_0_wdata2 : reg_type5_data_3_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_179 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h11 ? reg_type5_data_3_2 : reg_type5_data_3_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_180 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h11 ? io_exe_wb_1_wdata1 : _GEN_176; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_181 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h11 ? reg_type5_data_3_0 : _GEN_177; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_182 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h11 ? io_exe_wb_1_wdata2 : _GEN_178; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_183 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h11 ? reg_type5_data_3_2 : _GEN_179; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_184 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11 ? io_exe_wb_2_wdata1 : _GEN_180; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_185 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11 ? reg_type5_data_3_0 : _GEN_181; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_186 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11 ? io_exe_wb_2_wdata2 : _GEN_182; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_187 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11 ? reg_type5_data_3_2 : _GEN_183; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_188 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11 ? io_exe_wb_3_wdata1 : _GEN_184; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_189 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11 ? reg_type5_data_3_0 : _GEN_185; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_190 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11 ? io_exe_wb_3_wdata2 : _GEN_186; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_191 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11 ? reg_type5_data_3_2 : _GEN_187; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_192 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11 ? io_exe_wb_4_wdata1 : _GEN_188; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_193 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11 ? reg_type5_data_3_0 : _GEN_189; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_194 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11 ? io_exe_wb_4_wdata2 : _GEN_190; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_195 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11 ? reg_type5_data_3_2 : _GEN_191; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_3_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11 ? 32'h0 : _GEN_192; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_3_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11 ? reg_type5_data_3_0 : _GEN_193; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_3_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11 ? io_exe_wb_5_wdata2 : _GEN_194; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_3_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11 ? reg_type5_data_3_2 : _GEN_195; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_4_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_4_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_4_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_4_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_200 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h12 ? io_exe_wb_0_wdata1 : reg_type5_data_4_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_201 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h12 ? reg_type5_data_4_0 : reg_type5_data_4_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_202 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h12 ? io_exe_wb_0_wdata2 : reg_type5_data_4_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_203 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h12 ? reg_type5_data_4_2 : reg_type5_data_4_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_204 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h12 ? io_exe_wb_1_wdata1 : _GEN_200; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_205 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h12 ? reg_type5_data_4_0 : _GEN_201; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_206 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h12 ? io_exe_wb_1_wdata2 : _GEN_202; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_207 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h12 ? reg_type5_data_4_2 : _GEN_203; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_208 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12 ? io_exe_wb_2_wdata1 : _GEN_204; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_209 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12 ? reg_type5_data_4_0 : _GEN_205; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_210 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12 ? io_exe_wb_2_wdata2 : _GEN_206; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_211 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12 ? reg_type5_data_4_2 : _GEN_207; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_212 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12 ? io_exe_wb_3_wdata1 : _GEN_208; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_213 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12 ? reg_type5_data_4_0 : _GEN_209; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_214 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12 ? io_exe_wb_3_wdata2 : _GEN_210; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_215 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12 ? reg_type5_data_4_2 : _GEN_211; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_216 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12 ? io_exe_wb_4_wdata1 : _GEN_212; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_217 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12 ? reg_type5_data_4_0 : _GEN_213; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_218 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12 ? io_exe_wb_4_wdata2 : _GEN_214; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_219 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12 ? reg_type5_data_4_2 : _GEN_215; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_4_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12 ? 32'h0 : _GEN_216; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_4_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12 ? reg_type5_data_4_0 : _GEN_217; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_4_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12 ? io_exe_wb_5_wdata2 : _GEN_218; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_4_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12 ? reg_type5_data_4_2 : _GEN_219; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_5_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_5_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_5_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_5_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_224 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h13 ? io_exe_wb_0_wdata1 : reg_type5_data_5_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_225 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h13 ? reg_type5_data_5_0 : reg_type5_data_5_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_226 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h13 ? io_exe_wb_0_wdata2 : reg_type5_data_5_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_227 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h13 ? reg_type5_data_5_2 : reg_type5_data_5_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_228 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h13 ? io_exe_wb_1_wdata1 : _GEN_224; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_229 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h13 ? reg_type5_data_5_0 : _GEN_225; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_230 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h13 ? io_exe_wb_1_wdata2 : _GEN_226; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_231 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h13 ? reg_type5_data_5_2 : _GEN_227; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_232 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13 ? io_exe_wb_2_wdata1 : _GEN_228; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_233 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13 ? reg_type5_data_5_0 : _GEN_229; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_234 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13 ? io_exe_wb_2_wdata2 : _GEN_230; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_235 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13 ? reg_type5_data_5_2 : _GEN_231; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_236 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13 ? io_exe_wb_3_wdata1 : _GEN_232; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_237 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13 ? reg_type5_data_5_0 : _GEN_233; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_238 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13 ? io_exe_wb_3_wdata2 : _GEN_234; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_239 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13 ? reg_type5_data_5_2 : _GEN_235; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_240 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13 ? io_exe_wb_4_wdata1 : _GEN_236; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_241 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13 ? reg_type5_data_5_0 : _GEN_237; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_242 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13 ? io_exe_wb_4_wdata2 : _GEN_238; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_243 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13 ? reg_type5_data_5_2 : _GEN_239; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_5_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13 ? 32'h0 : _GEN_240; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_5_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13 ? reg_type5_data_5_0 : _GEN_241; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_5_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13 ? io_exe_wb_5_wdata2 : _GEN_242; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_5_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13 ? reg_type5_data_5_2 : _GEN_243; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_6_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_6_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_6_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_6_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_248 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h14 ? io_exe_wb_0_wdata1 : reg_type5_data_6_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_249 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h14 ? reg_type5_data_6_0 : reg_type5_data_6_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_250 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h14 ? io_exe_wb_0_wdata2 : reg_type5_data_6_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_251 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h14 ? reg_type5_data_6_2 : reg_type5_data_6_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_252 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h14 ? io_exe_wb_1_wdata1 : _GEN_248; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_253 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h14 ? reg_type5_data_6_0 : _GEN_249; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_254 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h14 ? io_exe_wb_1_wdata2 : _GEN_250; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_255 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h14 ? reg_type5_data_6_2 : _GEN_251; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_256 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14 ? io_exe_wb_2_wdata1 : _GEN_252; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_257 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14 ? reg_type5_data_6_0 : _GEN_253; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_258 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14 ? io_exe_wb_2_wdata2 : _GEN_254; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_259 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14 ? reg_type5_data_6_2 : _GEN_255; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_260 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14 ? io_exe_wb_3_wdata1 : _GEN_256; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_261 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14 ? reg_type5_data_6_0 : _GEN_257; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_262 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14 ? io_exe_wb_3_wdata2 : _GEN_258; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_263 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14 ? reg_type5_data_6_2 : _GEN_259; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_264 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14 ? io_exe_wb_4_wdata1 : _GEN_260; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_265 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14 ? reg_type5_data_6_0 : _GEN_261; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_266 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14 ? io_exe_wb_4_wdata2 : _GEN_262; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_267 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14 ? reg_type5_data_6_2 : _GEN_263; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_6_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14 ? 32'h0 : _GEN_264; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_6_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14 ? reg_type5_data_6_0 : _GEN_265; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_6_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14 ? io_exe_wb_5_wdata2 : _GEN_266; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_6_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14 ? reg_type5_data_6_2 : _GEN_267; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_7_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_7_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_7_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_7_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_272 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h15 ? io_exe_wb_0_wdata1 : reg_type5_data_7_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_273 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h15 ? reg_type5_data_7_0 : reg_type5_data_7_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_274 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h15 ? io_exe_wb_0_wdata2 : reg_type5_data_7_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_275 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h15 ? reg_type5_data_7_2 : reg_type5_data_7_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_276 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h15 ? io_exe_wb_1_wdata1 : _GEN_272; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_277 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h15 ? reg_type5_data_7_0 : _GEN_273; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_278 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h15 ? io_exe_wb_1_wdata2 : _GEN_274; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_279 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h15 ? reg_type5_data_7_2 : _GEN_275; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_280 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15 ? io_exe_wb_2_wdata1 : _GEN_276; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_281 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15 ? reg_type5_data_7_0 : _GEN_277; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_282 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15 ? io_exe_wb_2_wdata2 : _GEN_278; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_283 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15 ? reg_type5_data_7_2 : _GEN_279; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_284 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15 ? io_exe_wb_3_wdata1 : _GEN_280; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_285 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15 ? reg_type5_data_7_0 : _GEN_281; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_286 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15 ? io_exe_wb_3_wdata2 : _GEN_282; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_287 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15 ? reg_type5_data_7_2 : _GEN_283; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_288 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15 ? io_exe_wb_4_wdata1 : _GEN_284; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_289 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15 ? reg_type5_data_7_0 : _GEN_285; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_290 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15 ? io_exe_wb_4_wdata2 : _GEN_286; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_291 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15 ? reg_type5_data_7_2 : _GEN_287; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_7_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15 ? 32'h0 : _GEN_288; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_7_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15 ? reg_type5_data_7_0 : _GEN_289; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_7_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15 ? io_exe_wb_5_wdata2 : _GEN_290; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_7_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15 ? reg_type5_data_7_2 : _GEN_291; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_8_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_8_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_8_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_8_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_296 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h16 ? io_exe_wb_0_wdata1 : reg_type5_data_8_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_297 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h16 ? reg_type5_data_8_0 : reg_type5_data_8_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_298 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h16 ? io_exe_wb_0_wdata2 : reg_type5_data_8_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_299 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h16 ? reg_type5_data_8_2 : reg_type5_data_8_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_300 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h16 ? io_exe_wb_1_wdata1 : _GEN_296; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_301 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h16 ? reg_type5_data_8_0 : _GEN_297; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_302 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h16 ? io_exe_wb_1_wdata2 : _GEN_298; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_303 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h16 ? reg_type5_data_8_2 : _GEN_299; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_304 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16 ? io_exe_wb_2_wdata1 : _GEN_300; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_305 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16 ? reg_type5_data_8_0 : _GEN_301; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_306 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16 ? io_exe_wb_2_wdata2 : _GEN_302; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_307 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16 ? reg_type5_data_8_2 : _GEN_303; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_308 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16 ? io_exe_wb_3_wdata1 : _GEN_304; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_309 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16 ? reg_type5_data_8_0 : _GEN_305; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_310 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16 ? io_exe_wb_3_wdata2 : _GEN_306; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_311 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16 ? reg_type5_data_8_2 : _GEN_307; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_312 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16 ? io_exe_wb_4_wdata1 : _GEN_308; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_313 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16 ? reg_type5_data_8_0 : _GEN_309; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_314 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16 ? io_exe_wb_4_wdata2 : _GEN_310; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_315 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16 ? reg_type5_data_8_2 : _GEN_311; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_8_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16 ? 32'h0 : _GEN_312; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_8_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16 ? reg_type5_data_8_0 : _GEN_313; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_8_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16 ? io_exe_wb_5_wdata2 : _GEN_314; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_8_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16 ? reg_type5_data_8_2 : _GEN_315; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_9_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_9_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_9_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_9_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_320 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h17 ? io_exe_wb_0_wdata1 : reg_type5_data_9_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_321 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h17 ? reg_type5_data_9_0 : reg_type5_data_9_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_322 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h17 ? io_exe_wb_0_wdata2 : reg_type5_data_9_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_323 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h17 ? reg_type5_data_9_2 : reg_type5_data_9_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_324 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h17 ? io_exe_wb_1_wdata1 : _GEN_320; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_325 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h17 ? reg_type5_data_9_0 : _GEN_321; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_326 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h17 ? io_exe_wb_1_wdata2 : _GEN_322; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_327 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h17 ? reg_type5_data_9_2 : _GEN_323; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_328 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17 ? io_exe_wb_2_wdata1 : _GEN_324; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_329 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17 ? reg_type5_data_9_0 : _GEN_325; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_330 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17 ? io_exe_wb_2_wdata2 : _GEN_326; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_331 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17 ? reg_type5_data_9_2 : _GEN_327; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_332 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17 ? io_exe_wb_3_wdata1 : _GEN_328; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_333 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17 ? reg_type5_data_9_0 : _GEN_329; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_334 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17 ? io_exe_wb_3_wdata2 : _GEN_330; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_335 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17 ? reg_type5_data_9_2 : _GEN_331; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_336 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17 ? io_exe_wb_4_wdata1 : _GEN_332; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_337 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17 ? reg_type5_data_9_0 : _GEN_333; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_338 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17 ? io_exe_wb_4_wdata2 : _GEN_334; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_339 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17 ? reg_type5_data_9_2 : _GEN_335; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_9_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17 ? 32'h0 : _GEN_336; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_9_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17 ? reg_type5_data_9_0 : _GEN_337; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_9_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17 ? io_exe_wb_5_wdata2 : _GEN_338; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_9_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17 ? reg_type5_data_9_2 : _GEN_339; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_10_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_10_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_10_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_10_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_344 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h18 ? io_exe_wb_0_wdata1 : reg_type5_data_10_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_345 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h18 ? reg_type5_data_10_0 : reg_type5_data_10_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_346 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h18 ? io_exe_wb_0_wdata2 : reg_type5_data_10_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_347 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h18 ? reg_type5_data_10_2 : reg_type5_data_10_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_348 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h18 ? io_exe_wb_1_wdata1 : _GEN_344; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_349 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h18 ? reg_type5_data_10_0 : _GEN_345; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_350 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h18 ? io_exe_wb_1_wdata2 : _GEN_346; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_351 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h18 ? reg_type5_data_10_2 : _GEN_347; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_352 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18 ? io_exe_wb_2_wdata1 : _GEN_348; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_353 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18 ? reg_type5_data_10_0 : _GEN_349; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_354 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18 ? io_exe_wb_2_wdata2 : _GEN_350; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_355 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18 ? reg_type5_data_10_2 : _GEN_351; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_356 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18 ? io_exe_wb_3_wdata1 : _GEN_352; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_357 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18 ? reg_type5_data_10_0 : _GEN_353; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_358 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18 ? io_exe_wb_3_wdata2 : _GEN_354; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_359 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18 ? reg_type5_data_10_2 : _GEN_355; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_360 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18 ? io_exe_wb_4_wdata1 : _GEN_356; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_361 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18 ? reg_type5_data_10_0 : _GEN_357; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_362 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18 ? io_exe_wb_4_wdata2 : _GEN_358; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_363 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18 ? reg_type5_data_10_2 : _GEN_359; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_10_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18 ? 32'h0 : _GEN_360; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_10_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18 ? reg_type5_data_10_0 : _GEN_361; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_10_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18 ? io_exe_wb_5_wdata2 : _GEN_362; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_10_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18 ? reg_type5_data_10_2 : _GEN_363; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_11_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_11_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_11_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_11_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_368 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h19 ? io_exe_wb_0_wdata1 : reg_type5_data_11_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_369 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h19 ? reg_type5_data_11_0 : reg_type5_data_11_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_370 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h19 ? io_exe_wb_0_wdata2 : reg_type5_data_11_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_371 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h19 ? reg_type5_data_11_2 : reg_type5_data_11_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_372 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h19 ? io_exe_wb_1_wdata1 : _GEN_368; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_373 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h19 ? reg_type5_data_11_0 : _GEN_369; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_374 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h19 ? io_exe_wb_1_wdata2 : _GEN_370; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_375 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h19 ? reg_type5_data_11_2 : _GEN_371; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_376 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19 ? io_exe_wb_2_wdata1 : _GEN_372; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_377 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19 ? reg_type5_data_11_0 : _GEN_373; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_378 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19 ? io_exe_wb_2_wdata2 : _GEN_374; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_379 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19 ? reg_type5_data_11_2 : _GEN_375; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_380 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19 ? io_exe_wb_3_wdata1 : _GEN_376; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_381 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19 ? reg_type5_data_11_0 : _GEN_377; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_382 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19 ? io_exe_wb_3_wdata2 : _GEN_378; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_383 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19 ? reg_type5_data_11_2 : _GEN_379; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_384 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19 ? io_exe_wb_4_wdata1 : _GEN_380; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_385 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19 ? reg_type5_data_11_0 : _GEN_381; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_386 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19 ? io_exe_wb_4_wdata2 : _GEN_382; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_387 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19 ? reg_type5_data_11_2 : _GEN_383; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_11_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19 ? 32'h0 : _GEN_384; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_11_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19 ? reg_type5_data_11_0 : _GEN_385; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_11_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19 ? io_exe_wb_5_wdata2 : _GEN_386; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_11_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19 ? reg_type5_data_11_2 : _GEN_387; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_12_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_12_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_12_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_12_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_392 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1a ? io_exe_wb_0_wdata1 : reg_type5_data_12_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_393 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1a ? reg_type5_data_12_0 : reg_type5_data_12_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_394 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1a ? io_exe_wb_0_wdata2 : reg_type5_data_12_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_395 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1a ? reg_type5_data_12_2 : reg_type5_data_12_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_396 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1a ? io_exe_wb_1_wdata1 : _GEN_392; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_397 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1a ? reg_type5_data_12_0 : _GEN_393; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_398 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1a ? io_exe_wb_1_wdata2 : _GEN_394; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_399 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1a ? reg_type5_data_12_2 : _GEN_395; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_400 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a ? io_exe_wb_2_wdata1 : _GEN_396; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_401 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a ? reg_type5_data_12_0 : _GEN_397; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_402 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a ? io_exe_wb_2_wdata2 : _GEN_398; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_403 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a ? reg_type5_data_12_2 : _GEN_399; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_404 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a ? io_exe_wb_3_wdata1 : _GEN_400; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_405 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a ? reg_type5_data_12_0 : _GEN_401; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_406 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a ? io_exe_wb_3_wdata2 : _GEN_402; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_407 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a ? reg_type5_data_12_2 : _GEN_403; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_408 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a ? io_exe_wb_4_wdata1 : _GEN_404; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_409 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a ? reg_type5_data_12_0 : _GEN_405; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_410 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a ? io_exe_wb_4_wdata2 : _GEN_406; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_411 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a ? reg_type5_data_12_2 : _GEN_407; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_12_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a ? 32'h0 : _GEN_408; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_12_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a ? reg_type5_data_12_0 : _GEN_409; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_12_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a ? io_exe_wb_5_wdata2 : _GEN_410; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_12_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a ? reg_type5_data_12_2 : _GEN_411; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_13_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_13_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_13_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_13_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_416 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1b ? io_exe_wb_0_wdata1 : reg_type5_data_13_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_417 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1b ? reg_type5_data_13_0 : reg_type5_data_13_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_418 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1b ? io_exe_wb_0_wdata2 : reg_type5_data_13_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_419 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1b ? reg_type5_data_13_2 : reg_type5_data_13_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_420 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1b ? io_exe_wb_1_wdata1 : _GEN_416; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_421 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1b ? reg_type5_data_13_0 : _GEN_417; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_422 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1b ? io_exe_wb_1_wdata2 : _GEN_418; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_423 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1b ? reg_type5_data_13_2 : _GEN_419; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_424 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b ? io_exe_wb_2_wdata1 : _GEN_420; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_425 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b ? reg_type5_data_13_0 : _GEN_421; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_426 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b ? io_exe_wb_2_wdata2 : _GEN_422; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_427 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b ? reg_type5_data_13_2 : _GEN_423; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_428 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b ? io_exe_wb_3_wdata1 : _GEN_424; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_429 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b ? reg_type5_data_13_0 : _GEN_425; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_430 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b ? io_exe_wb_3_wdata2 : _GEN_426; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_431 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b ? reg_type5_data_13_2 : _GEN_427; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_432 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b ? io_exe_wb_4_wdata1 : _GEN_428; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_433 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b ? reg_type5_data_13_0 : _GEN_429; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_434 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b ? io_exe_wb_4_wdata2 : _GEN_430; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_435 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b ? reg_type5_data_13_2 : _GEN_431; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_13_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b ? 32'h0 : _GEN_432; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_13_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b ? reg_type5_data_13_0 : _GEN_433; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_13_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b ? io_exe_wb_5_wdata2 : _GEN_434; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_13_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b ? reg_type5_data_13_2 : _GEN_435; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_14_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_14_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_14_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_14_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_440 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1c ? io_exe_wb_0_wdata1 : reg_type5_data_14_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_441 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1c ? reg_type5_data_14_0 : reg_type5_data_14_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_442 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1c ? io_exe_wb_0_wdata2 : reg_type5_data_14_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_443 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1c ? reg_type5_data_14_2 : reg_type5_data_14_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_444 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1c ? io_exe_wb_1_wdata1 : _GEN_440; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_445 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1c ? reg_type5_data_14_0 : _GEN_441; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_446 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1c ? io_exe_wb_1_wdata2 : _GEN_442; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_447 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1c ? reg_type5_data_14_2 : _GEN_443; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_448 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c ? io_exe_wb_2_wdata1 : _GEN_444; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_449 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c ? reg_type5_data_14_0 : _GEN_445; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_450 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c ? io_exe_wb_2_wdata2 : _GEN_446; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_451 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c ? reg_type5_data_14_2 : _GEN_447; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_452 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c ? io_exe_wb_3_wdata1 : _GEN_448; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_453 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c ? reg_type5_data_14_0 : _GEN_449; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_454 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c ? io_exe_wb_3_wdata2 : _GEN_450; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_455 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c ? reg_type5_data_14_2 : _GEN_451; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_456 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c ? io_exe_wb_4_wdata1 : _GEN_452; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_457 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c ? reg_type5_data_14_0 : _GEN_453; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_458 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c ? io_exe_wb_4_wdata2 : _GEN_454; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_459 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c ? reg_type5_data_14_2 : _GEN_455; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_14_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c ? 32'h0 : _GEN_456; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_14_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c ? reg_type5_data_14_0 : _GEN_457; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_14_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c ? io_exe_wb_5_wdata2 : _GEN_458; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_14_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c ? reg_type5_data_14_2 : _GEN_459; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_15_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_15_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_15_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_15_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_464 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1d ? io_exe_wb_0_wdata1 : reg_type5_data_15_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_465 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1d ? reg_type5_data_15_0 : reg_type5_data_15_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_466 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1d ? io_exe_wb_0_wdata2 : reg_type5_data_15_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_467 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1d ? reg_type5_data_15_2 : reg_type5_data_15_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_468 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1d ? io_exe_wb_1_wdata1 : _GEN_464; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_469 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1d ? reg_type5_data_15_0 : _GEN_465; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_470 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1d ? io_exe_wb_1_wdata2 : _GEN_466; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_471 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1d ? reg_type5_data_15_2 : _GEN_467; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_472 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d ? io_exe_wb_2_wdata1 : _GEN_468; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_473 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d ? reg_type5_data_15_0 : _GEN_469; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_474 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d ? io_exe_wb_2_wdata2 : _GEN_470; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_475 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d ? reg_type5_data_15_2 : _GEN_471; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_476 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d ? io_exe_wb_3_wdata1 : _GEN_472; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_477 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d ? reg_type5_data_15_0 : _GEN_473; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_478 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d ? io_exe_wb_3_wdata2 : _GEN_474; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_479 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d ? reg_type5_data_15_2 : _GEN_475; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_480 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d ? io_exe_wb_4_wdata1 : _GEN_476; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_481 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d ? reg_type5_data_15_0 : _GEN_477; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_482 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d ? io_exe_wb_4_wdata2 : _GEN_478; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_483 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d ? reg_type5_data_15_2 : _GEN_479; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_15_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d ? 32'h0 : _GEN_480; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_15_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d ? reg_type5_data_15_0 : _GEN_481; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_15_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d ? io_exe_wb_5_wdata2 : _GEN_482; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_15_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d ? reg_type5_data_15_2 : _GEN_483; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_16_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_16_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_16_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_16_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_488 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1e ? io_exe_wb_0_wdata1 : reg_type5_data_16_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_489 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1e ? reg_type5_data_16_0 : reg_type5_data_16_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_490 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1e ? io_exe_wb_0_wdata2 : reg_type5_data_16_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_491 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1e ? reg_type5_data_16_2 : reg_type5_data_16_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_492 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1e ? io_exe_wb_1_wdata1 : _GEN_488; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_493 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1e ? reg_type5_data_16_0 : _GEN_489; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_494 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1e ? io_exe_wb_1_wdata2 : _GEN_490; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_495 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1e ? reg_type5_data_16_2 : _GEN_491; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_496 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e ? io_exe_wb_2_wdata1 : _GEN_492; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_497 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e ? reg_type5_data_16_0 : _GEN_493; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_498 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e ? io_exe_wb_2_wdata2 : _GEN_494; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_499 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e ? reg_type5_data_16_2 : _GEN_495; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_500 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e ? io_exe_wb_3_wdata1 : _GEN_496; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_501 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e ? reg_type5_data_16_0 : _GEN_497; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_502 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e ? io_exe_wb_3_wdata2 : _GEN_498; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_503 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e ? reg_type5_data_16_2 : _GEN_499; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_504 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e ? io_exe_wb_4_wdata1 : _GEN_500; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_505 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e ? reg_type5_data_16_0 : _GEN_501; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_506 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e ? io_exe_wb_4_wdata2 : _GEN_502; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_507 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e ? reg_type5_data_16_2 : _GEN_503; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_16_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e ? 32'h0 : _GEN_504; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_16_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e ? reg_type5_data_16_0 : _GEN_505; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_16_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e ? io_exe_wb_5_wdata2 : _GEN_506; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_16_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e ? reg_type5_data_16_2 : _GEN_507; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_17_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_17_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_17_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_17_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_512 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1f ? io_exe_wb_0_wdata1 : reg_type5_data_17_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_513 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1f ? reg_type5_data_17_0 : reg_type5_data_17_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_514 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1f ? io_exe_wb_0_wdata2 : reg_type5_data_17_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_515 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h1f ? reg_type5_data_17_2 : reg_type5_data_17_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_516 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1f ? io_exe_wb_1_wdata1 : _GEN_512; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_517 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1f ? reg_type5_data_17_0 : _GEN_513; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_518 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1f ? io_exe_wb_1_wdata2 : _GEN_514; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_519 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h1f ? reg_type5_data_17_2 : _GEN_515; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_520 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f ? io_exe_wb_2_wdata1 : _GEN_516; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_521 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f ? reg_type5_data_17_0 : _GEN_517; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_522 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f ? io_exe_wb_2_wdata2 : _GEN_518; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_523 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f ? reg_type5_data_17_2 : _GEN_519; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_524 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f ? io_exe_wb_3_wdata1 : _GEN_520; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_525 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f ? reg_type5_data_17_0 : _GEN_521; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_526 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f ? io_exe_wb_3_wdata2 : _GEN_522; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_527 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f ? reg_type5_data_17_2 : _GEN_523; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_528 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f ? io_exe_wb_4_wdata1 : _GEN_524; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_529 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f ? reg_type5_data_17_0 : _GEN_525; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_530 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f ? io_exe_wb_4_wdata2 : _GEN_526; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_531 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f ? reg_type5_data_17_2 : _GEN_527; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_17_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f ? 32'h0 : _GEN_528; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_17_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f ? reg_type5_data_17_0 : _GEN_529; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_17_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f ? io_exe_wb_5_wdata2 : _GEN_530; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_17_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f ? reg_type5_data_17_2 : _GEN_531; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_18_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_18_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_18_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_18_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_536 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h20 ? io_exe_wb_0_wdata1 : reg_type5_data_18_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_537 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h20 ? reg_type5_data_18_0 : reg_type5_data_18_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_538 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h20 ? io_exe_wb_0_wdata2 : reg_type5_data_18_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_539 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h20 ? reg_type5_data_18_2 : reg_type5_data_18_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_540 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h20 ? io_exe_wb_1_wdata1 : _GEN_536; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_541 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h20 ? reg_type5_data_18_0 : _GEN_537; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_542 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h20 ? io_exe_wb_1_wdata2 : _GEN_538; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_543 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h20 ? reg_type5_data_18_2 : _GEN_539; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_544 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20 ? io_exe_wb_2_wdata1 : _GEN_540; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_545 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20 ? reg_type5_data_18_0 : _GEN_541; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_546 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20 ? io_exe_wb_2_wdata2 : _GEN_542; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_547 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20 ? reg_type5_data_18_2 : _GEN_543; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_548 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20 ? io_exe_wb_3_wdata1 : _GEN_544; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_549 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20 ? reg_type5_data_18_0 : _GEN_545; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_550 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20 ? io_exe_wb_3_wdata2 : _GEN_546; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_551 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20 ? reg_type5_data_18_2 : _GEN_547; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_552 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20 ? io_exe_wb_4_wdata1 : _GEN_548; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_553 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20 ? reg_type5_data_18_0 : _GEN_549; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_554 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20 ? io_exe_wb_4_wdata2 : _GEN_550; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_555 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20 ? reg_type5_data_18_2 : _GEN_551; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_18_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20 ? 32'h0 : _GEN_552; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_18_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20 ? reg_type5_data_18_0 : _GEN_553; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_18_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20 ? io_exe_wb_5_wdata2 : _GEN_554; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_18_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20 ? reg_type5_data_18_2 : _GEN_555; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_19_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_19_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_19_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_19_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_560 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h21 ? io_exe_wb_0_wdata1 : reg_type5_data_19_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_561 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h21 ? reg_type5_data_19_0 : reg_type5_data_19_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_562 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h21 ? io_exe_wb_0_wdata2 : reg_type5_data_19_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_563 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h21 ? reg_type5_data_19_2 : reg_type5_data_19_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_564 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h21 ? io_exe_wb_1_wdata1 : _GEN_560; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_565 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h21 ? reg_type5_data_19_0 : _GEN_561; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_566 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h21 ? io_exe_wb_1_wdata2 : _GEN_562; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_567 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h21 ? reg_type5_data_19_2 : _GEN_563; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_568 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21 ? io_exe_wb_2_wdata1 : _GEN_564; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_569 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21 ? reg_type5_data_19_0 : _GEN_565; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_570 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21 ? io_exe_wb_2_wdata2 : _GEN_566; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_571 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21 ? reg_type5_data_19_2 : _GEN_567; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_572 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21 ? io_exe_wb_3_wdata1 : _GEN_568; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_573 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21 ? reg_type5_data_19_0 : _GEN_569; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_574 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21 ? io_exe_wb_3_wdata2 : _GEN_570; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_575 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21 ? reg_type5_data_19_2 : _GEN_571; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_576 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21 ? io_exe_wb_4_wdata1 : _GEN_572; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_577 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21 ? reg_type5_data_19_0 : _GEN_573; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_578 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21 ? io_exe_wb_4_wdata2 : _GEN_574; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_579 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21 ? reg_type5_data_19_2 : _GEN_575; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_19_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21 ? 32'h0 : _GEN_576; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_19_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21 ? reg_type5_data_19_0 : _GEN_577; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_19_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21 ? io_exe_wb_5_wdata2 : _GEN_578; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_19_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21 ? reg_type5_data_19_2 : _GEN_579; // @[regfile.scala 51:64 regfile.scala 56:27]
  reg [31:0] reg_type5_data_20_0; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_20_1; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_20_2; // @[regfile.scala 22:22]
  reg [31:0] reg_type5_data_20_3; // @[regfile.scala 22:22]
  wire [31:0] _GEN_584 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h22 ? io_exe_wb_0_wdata1 : reg_type5_data_20_0; // @[regfile.scala 51:64 regfile.scala 53:27 regfile.scala 40:18]
  wire [31:0] _GEN_585 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h22 ? reg_type5_data_20_0 : reg_type5_data_20_1; // @[regfile.scala 51:64 regfile.scala 54:27 regfile.scala 40:18]
  wire [31:0] _GEN_586 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h22 ? io_exe_wb_0_wdata2 : reg_type5_data_20_2; // @[regfile.scala 51:64 regfile.scala 55:27 regfile.scala 40:18]
  wire [31:0] _GEN_587 = io_exe_wb_0_vld & io_exe_wb_0_gregidx == 6'h22 ? reg_type5_data_20_2 : reg_type5_data_20_3; // @[regfile.scala 51:64 regfile.scala 56:27 regfile.scala 40:18]
  wire [31:0] _GEN_588 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h22 ? io_exe_wb_1_wdata1 : _GEN_584; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_589 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h22 ? reg_type5_data_20_0 : _GEN_585; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_590 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h22 ? io_exe_wb_1_wdata2 : _GEN_586; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_591 = io_exe_wb_1_vld & io_exe_wb_1_gregidx == 6'h22 ? reg_type5_data_20_2 : _GEN_587; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_592 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22 ? io_exe_wb_2_wdata1 : _GEN_588; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_593 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22 ? reg_type5_data_20_0 : _GEN_589; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_594 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22 ? io_exe_wb_2_wdata2 : _GEN_590; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_595 = io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22 ? reg_type5_data_20_2 : _GEN_591; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_596 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22 ? io_exe_wb_3_wdata1 : _GEN_592; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_597 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22 ? reg_type5_data_20_0 : _GEN_593; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_598 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22 ? io_exe_wb_3_wdata2 : _GEN_594; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_599 = io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22 ? reg_type5_data_20_2 : _GEN_595; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] _GEN_600 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22 ? io_exe_wb_4_wdata1 : _GEN_596; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] _GEN_601 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22 ? reg_type5_data_20_0 : _GEN_597; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] _GEN_602 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22 ? io_exe_wb_4_wdata2 : _GEN_598; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] _GEN_603 = io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22 ? reg_type5_data_20_2 : _GEN_599; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] reg_type5_data_nxt_20_0 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22 ? 32'h0 : _GEN_600; // @[regfile.scala 51:64 regfile.scala 53:27]
  wire [31:0] reg_type5_data_nxt_20_1 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22 ? reg_type5_data_20_0 : _GEN_601; // @[regfile.scala 51:64 regfile.scala 54:27]
  wire [31:0] reg_type5_data_nxt_20_2 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22 ? io_exe_wb_5_wdata2 : _GEN_602; // @[regfile.scala 51:64 regfile.scala 55:27]
  wire [31:0] reg_type5_data_nxt_20_3 = io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22 ? reg_type5_data_20_2 : _GEN_603; // @[regfile.scala 51:64 regfile.scala 56:27]
  wire [31:0] tmp_0_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out = io_exe_rd_0_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_617 = io_exe_rd_0_req_gidx[0] ? io_coef_in_mainch_drc_smooth_1 : io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out = io_exe_rd_0_req_gidx < 3'h2 ? _GEN_617 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out = io_exe_rd_0_req_iscoef ? tmp_8_out_out_out : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_621 = io_exe_rd_0_req_gidx[0] ? io_coef_in_subch_drc_smooth_1 : io_coef_in_subch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out = io_exe_rd_0_req_gidx < 3'h2 ? _GEN_621 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out = io_exe_rd_0_req_iscoef ? tmp_9_out_out_out : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_625 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_626 = 3'h2 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_625; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_627 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_626; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_628 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_627; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_628 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out = io_exe_rd_0_req_iscoef ? tmp_10_out_out_out : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out = io_exe_rd_0_req_iscoef ? tmp_10_out_out_out : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_639 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_640 = 3'h2 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_639; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_641 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_640; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_642 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_641; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_642 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out = io_exe_rd_0_req_iscoef ? tmp_12_out_out_out : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out = io_exe_rd_0_req_iscoef ? tmp_12_out_out_out : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_653 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_654 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_653; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_655 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_654; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_656 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_655; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_656 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_2 = io_exe_rd_0_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_659 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_660 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt__2 : _GEN_659; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_661 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt__3 : _GEN_660; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_661 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_14_out_out_out_1 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out = io_exe_rd_0_req_iscoef ? tmp_14_out_out_out : tmp_14_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_666 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_667 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_666; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_668 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_667; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_669 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_668; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_669 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_672 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_673 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_1_2 : _GEN_672; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_674 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_1_3 : _GEN_673; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_674 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_15_out_out_out_1 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out = io_exe_rd_0_req_iscoef ? tmp_15_out_out_out : tmp_15_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_679 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_680 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_679; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_681 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_680; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_682 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_681; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_682 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_685 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_686 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_2_2 : _GEN_685; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_687 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_2_3 : _GEN_686; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_687 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_16_out_out_out_1 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out = io_exe_rd_0_req_iscoef ? tmp_16_out_out_out : tmp_16_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_692 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_693 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_692; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_694 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_693; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_695 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_694; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_695 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_698 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_699 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_3_2 : _GEN_698; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_700 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_3_3 : _GEN_699; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_700 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_17_out_out_out_1 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out = io_exe_rd_0_req_iscoef ? tmp_17_out_out_out : tmp_17_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_705 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_706 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_705; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_707 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_706; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_708 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_707; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_708 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_711 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_712 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_4_2 : _GEN_711; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_713 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_4_3 : _GEN_712; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_713 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_18_out_out_out_1 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out = io_exe_rd_0_req_iscoef ? tmp_18_out_out_out : tmp_18_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_718 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_719 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_718; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_720 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_719; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_721 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_720; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_721 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_724 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_725 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_5_2 : _GEN_724; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_726 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_5_3 : _GEN_725; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_726 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_19_out_out_out_1 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out = io_exe_rd_0_req_iscoef ? tmp_19_out_out_out : tmp_19_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_731 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_732 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_731; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_733 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_732; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_734 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_733; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_734 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_737 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_738 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_6_2 : _GEN_737; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_739 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_6_3 : _GEN_738; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_739 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_20_out_out_out_1 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out = io_exe_rd_0_req_iscoef ? tmp_20_out_out_out : tmp_20_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_744 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_745 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_744; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_746 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_745; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_747 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_746; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_747 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_750 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_751 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_7_2 : _GEN_750; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_752 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_7_3 : _GEN_751; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_752 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_21_out_out_out_1 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out = io_exe_rd_0_req_iscoef ? tmp_21_out_out_out : tmp_21_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_757 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_758 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_757; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_759 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_758; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_760 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_759; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_760 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_763 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_764 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_8_2 : _GEN_763; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_765 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_8_3 : _GEN_764; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_765 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_22_out_out_out_1 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out = io_exe_rd_0_req_iscoef ? tmp_22_out_out_out : tmp_22_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_770 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_771 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_770; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_772 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_771; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_773 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_772; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_773 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_776 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_777 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_9_2 : _GEN_776; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_778 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_9_3 : _GEN_777; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_778 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_23_out_out_out_1 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out = io_exe_rd_0_req_iscoef ? tmp_23_out_out_out : tmp_23_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_783 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_784 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_783; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_785 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_784; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_786 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_785; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_786 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_789 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_790 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_10_2 : _GEN_789; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_791 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_10_3 : _GEN_790; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_791 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_24_out_out_out_1 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out = io_exe_rd_0_req_iscoef ? tmp_24_out_out_out : tmp_24_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_796 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_797 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_796; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_798 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_797; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_799 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_798; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_799 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_802 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_803 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_11_2 : _GEN_802; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_804 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_11_3 : _GEN_803; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_804 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_25_out_out_out_1 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out = io_exe_rd_0_req_iscoef ? tmp_25_out_out_out : tmp_25_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_809 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_810 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_809; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_811 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_810; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_812 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_811; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_812 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_815 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_816 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_12_2 : _GEN_815; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_817 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_12_3 : _GEN_816; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_817 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_26_out_out_out_1 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out = io_exe_rd_0_req_iscoef ? tmp_26_out_out_out : tmp_26_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_822 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_823 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_822; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_824 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_823; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_825 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_824; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_825 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_828 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_829 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_13_2 : _GEN_828; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_830 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_13_3 : _GEN_829; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_830 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_27_out_out_out_1 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out = io_exe_rd_0_req_iscoef ? tmp_27_out_out_out : tmp_27_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_835 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_836 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_835; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_837 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_836; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_838 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_837; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_838 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_841 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_842 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_14_2 : _GEN_841; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_843 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_14_3 : _GEN_842; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_843 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_28_out_out_out_1 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out = io_exe_rd_0_req_iscoef ? tmp_28_out_out_out : tmp_28_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_848 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_849 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_848; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_850 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_849; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_851 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_850; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_851 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_854 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_855 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_15_2 : _GEN_854; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_856 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_15_3 : _GEN_855; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_856 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_29_out_out_out_1 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out = io_exe_rd_0_req_iscoef ? tmp_29_out_out_out : tmp_29_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_861 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_862 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_861; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_863 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_862; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_864 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_863; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_864 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_867 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_868 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_16_2 : _GEN_867; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_869 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_16_3 : _GEN_868; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_869 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_30_out_out_out_1 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out = io_exe_rd_0_req_iscoef ? tmp_30_out_out_out : tmp_30_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_874 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_875 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_874; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_876 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_875; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_877 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_876; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_877 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_880 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_881 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_17_2 : _GEN_880; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_882 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_17_3 : _GEN_881; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_882 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_31_out_out_out_1 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out = io_exe_rd_0_req_iscoef ? tmp_31_out_out_out : tmp_31_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_887 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_888 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_887; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_889 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_888; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_890 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_889; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_890 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_893 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_894 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_18_2 : _GEN_893; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_895 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_18_3 : _GEN_894; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_895 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_32_out_out_out_1 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out = io_exe_rd_0_req_iscoef ? tmp_32_out_out_out : tmp_32_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_900 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_901 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_900; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_902 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_901; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_903 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_902; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_903 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_906 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_907 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_19_2 : _GEN_906; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_908 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_19_3 : _GEN_907; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_908 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_33_out_out_out_1 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out = io_exe_rd_0_req_iscoef ? tmp_33_out_out_out : tmp_33_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_913 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_914 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_913; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_915 = 3'h3 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_914; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_916 = 3'h4 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_915; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_916 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_919 = 2'h1 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_920 = 2'h2 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_20_2 : _GEN_919; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_921 = 2'h3 == _tmp_14_out_out_T_2[1:0] ? reg_type5_data_nxt_20_3 : _GEN_920; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_1 = _tmp_14_out_out_T_2 < 3'h4 ? _GEN_921 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_1 = io_exe_rd_0_req_isgroup ? tmp_34_out_out_out_1 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out = io_exe_rd_0_req_iscoef ? tmp_34_out_out_out : tmp_34_out_out_1; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_926 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_927 = 3'h2 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_926; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_928 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_927; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_929 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_928; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_929 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out = io_exe_rd_0_req_iscoef ? tmp_35_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_933 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_934 = 3'h2 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_933; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_935 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_934; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_936 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_935; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_936 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out = io_exe_rd_0_req_iscoef ? tmp_36_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_940 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_941 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_940; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_942 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_941; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_943 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_942; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_943 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out = io_exe_rd_0_req_iscoef ? tmp_37_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_947 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_948 = 3'h2 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_947; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_949 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_948; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_950 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_949; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_950 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out = io_exe_rd_0_req_iscoef ? tmp_38_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_954 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_955 = 3'h2 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_954; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_956 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_955; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_957 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_956; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_957 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out = io_exe_rd_0_req_iscoef ? tmp_39_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_961 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_962 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_961; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_963 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_962; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_964 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_963; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_964 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out = io_exe_rd_0_req_iscoef ? tmp_40_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_968 = 3'h1 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_969 = 3'h2 == io_exe_rd_0_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_968; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_970 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_969; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_971 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_970; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_971 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out = io_exe_rd_0_req_iscoef ? tmp_41_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] reg_type6_coef_7_0 = io_coef_in_subch_ch3sel ? 32'h0 : io_coef_in_subch_ch3mix_0; // @[regfile.scala 266:34]
  wire [31:0] reg_type6_coef_7_1 = io_coef_in_subch_ch3sel ? 32'h0 : io_coef_in_subch_ch3mix_1; // @[regfile.scala 267:34]
  wire [31:0] _GEN_975 = 3'h1 == io_exe_rd_0_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [23:0] _coef_2_T_1 = io_coef_in_subch_ch3sel ? 24'h800000 : 24'h0; // @[regfile.scala 268:34]
  wire [31:0] reg_type6_coef_7_2 = {{8'd0}, _coef_2_T_1}; // @[regfile.scala 24:38 regfile.scala 268:28]
  wire [31:0] _GEN_976 = 3'h2 == io_exe_rd_0_req_gidx ? reg_type6_coef_7_2 : _GEN_975; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_977 = 3'h3 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_976; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_978 = 3'h4 == io_exe_rd_0_req_gidx ? 32'h0 : _GEN_977; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out = io_exe_rd_0_req_gidx < 3'h5 ? _GEN_978 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out = io_exe_rd_0_req_iscoef ? tmp_42_out_out_out : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out = io_exe_rd_0_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out = io_exe_rd_0_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] reg_type7_coef_2_0 = io_coef_in_subch_ch2volsel ? io_coef_in_subch_ch2vol : io_coef_in_mainch_ch1_vol; // @[regfile.scala 272:34]
  wire [31:0] tmp_45_out = io_exe_rd_0_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] reg_type7_coef_3_0 = io_coef_in_subch_ch3volsel ? io_coef_in_subch_ch3vol : io_coef_in_mainch_ch0_vol; // @[regfile.scala 273:34]
  wire [31:0] tmp_46_out = io_exe_rd_0_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out = io_exe_rd_0_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out = io_exe_rd_0_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out = io_exe_rd_0_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out = io_exe_rd_0_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_0_resp_T = 64'h1 << io_exe_rd_0_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_0_resp_T_52 = _io_exe_rd_0_resp_T[0] ? tmp_0_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_53 = _io_exe_rd_0_resp_T[1] ? tmp_1_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_54 = _io_exe_rd_0_resp_T[2] ? tmp_2_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_55 = _io_exe_rd_0_resp_T[3] ? tmp_3_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_56 = _io_exe_rd_0_resp_T[4] ? tmp_4_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_57 = _io_exe_rd_0_resp_T[5] ? tmp_5_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_58 = _io_exe_rd_0_resp_T[6] ? tmp_6_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_59 = _io_exe_rd_0_resp_T[7] ? tmp_7_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_60 = _io_exe_rd_0_resp_T[8] ? tmp_8_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_61 = _io_exe_rd_0_resp_T[9] ? tmp_9_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_62 = _io_exe_rd_0_resp_T[10] ? tmp_10_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_63 = _io_exe_rd_0_resp_T[11] ? tmp_11_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_64 = _io_exe_rd_0_resp_T[12] ? tmp_12_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_65 = _io_exe_rd_0_resp_T[13] ? tmp_13_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_66 = _io_exe_rd_0_resp_T[14] ? tmp_14_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_67 = _io_exe_rd_0_resp_T[15] ? tmp_15_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_68 = _io_exe_rd_0_resp_T[16] ? tmp_16_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_69 = _io_exe_rd_0_resp_T[17] ? tmp_17_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_70 = _io_exe_rd_0_resp_T[18] ? tmp_18_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_71 = _io_exe_rd_0_resp_T[19] ? tmp_19_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_72 = _io_exe_rd_0_resp_T[20] ? tmp_20_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_73 = _io_exe_rd_0_resp_T[21] ? tmp_21_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_74 = _io_exe_rd_0_resp_T[22] ? tmp_22_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_75 = _io_exe_rd_0_resp_T[23] ? tmp_23_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_76 = _io_exe_rd_0_resp_T[24] ? tmp_24_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_77 = _io_exe_rd_0_resp_T[25] ? tmp_25_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_78 = _io_exe_rd_0_resp_T[26] ? tmp_26_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_79 = _io_exe_rd_0_resp_T[27] ? tmp_27_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_80 = _io_exe_rd_0_resp_T[28] ? tmp_28_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_81 = _io_exe_rd_0_resp_T[29] ? tmp_29_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_82 = _io_exe_rd_0_resp_T[30] ? tmp_30_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_83 = _io_exe_rd_0_resp_T[31] ? tmp_31_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_84 = _io_exe_rd_0_resp_T[32] ? tmp_32_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_85 = _io_exe_rd_0_resp_T[33] ? tmp_33_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_86 = _io_exe_rd_0_resp_T[34] ? tmp_34_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_87 = _io_exe_rd_0_resp_T[35] ? tmp_35_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_88 = _io_exe_rd_0_resp_T[36] ? tmp_36_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_89 = _io_exe_rd_0_resp_T[37] ? tmp_37_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_90 = _io_exe_rd_0_resp_T[38] ? tmp_38_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_91 = _io_exe_rd_0_resp_T[39] ? tmp_39_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_92 = _io_exe_rd_0_resp_T[40] ? tmp_40_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_93 = _io_exe_rd_0_resp_T[41] ? tmp_41_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_94 = _io_exe_rd_0_resp_T[42] ? tmp_42_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_95 = _io_exe_rd_0_resp_T[43] ? tmp_43_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_96 = _io_exe_rd_0_resp_T[44] ? tmp_44_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_97 = _io_exe_rd_0_resp_T[45] ? tmp_45_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_98 = _io_exe_rd_0_resp_T[46] ? tmp_46_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_99 = _io_exe_rd_0_resp_T[47] ? tmp_47_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_100 = _io_exe_rd_0_resp_T[48] ? tmp_48_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_101 = _io_exe_rd_0_resp_T[49] ? tmp_49_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_102 = _io_exe_rd_0_resp_T[50] ? tmp_50_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_103 = _io_exe_rd_0_resp_T_52 | _io_exe_rd_0_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_104 = _io_exe_rd_0_resp_T_103 | _io_exe_rd_0_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_105 = _io_exe_rd_0_resp_T_104 | _io_exe_rd_0_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_106 = _io_exe_rd_0_resp_T_105 | _io_exe_rd_0_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_107 = _io_exe_rd_0_resp_T_106 | _io_exe_rd_0_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_108 = _io_exe_rd_0_resp_T_107 | _io_exe_rd_0_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_109 = _io_exe_rd_0_resp_T_108 | _io_exe_rd_0_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_110 = _io_exe_rd_0_resp_T_109 | _io_exe_rd_0_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_111 = _io_exe_rd_0_resp_T_110 | _io_exe_rd_0_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_112 = _io_exe_rd_0_resp_T_111 | _io_exe_rd_0_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_113 = _io_exe_rd_0_resp_T_112 | _io_exe_rd_0_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_114 = _io_exe_rd_0_resp_T_113 | _io_exe_rd_0_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_115 = _io_exe_rd_0_resp_T_114 | _io_exe_rd_0_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_116 = _io_exe_rd_0_resp_T_115 | _io_exe_rd_0_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_117 = _io_exe_rd_0_resp_T_116 | _io_exe_rd_0_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_118 = _io_exe_rd_0_resp_T_117 | _io_exe_rd_0_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_119 = _io_exe_rd_0_resp_T_118 | _io_exe_rd_0_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_120 = _io_exe_rd_0_resp_T_119 | _io_exe_rd_0_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_121 = _io_exe_rd_0_resp_T_120 | _io_exe_rd_0_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_122 = _io_exe_rd_0_resp_T_121 | _io_exe_rd_0_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_123 = _io_exe_rd_0_resp_T_122 | _io_exe_rd_0_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_124 = _io_exe_rd_0_resp_T_123 | _io_exe_rd_0_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_125 = _io_exe_rd_0_resp_T_124 | _io_exe_rd_0_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_126 = _io_exe_rd_0_resp_T_125 | _io_exe_rd_0_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_127 = _io_exe_rd_0_resp_T_126 | _io_exe_rd_0_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_128 = _io_exe_rd_0_resp_T_127 | _io_exe_rd_0_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_129 = _io_exe_rd_0_resp_T_128 | _io_exe_rd_0_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_130 = _io_exe_rd_0_resp_T_129 | _io_exe_rd_0_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_131 = _io_exe_rd_0_resp_T_130 | _io_exe_rd_0_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_132 = _io_exe_rd_0_resp_T_131 | _io_exe_rd_0_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_133 = _io_exe_rd_0_resp_T_132 | _io_exe_rd_0_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_134 = _io_exe_rd_0_resp_T_133 | _io_exe_rd_0_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_135 = _io_exe_rd_0_resp_T_134 | _io_exe_rd_0_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_136 = _io_exe_rd_0_resp_T_135 | _io_exe_rd_0_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_137 = _io_exe_rd_0_resp_T_136 | _io_exe_rd_0_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_138 = _io_exe_rd_0_resp_T_137 | _io_exe_rd_0_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_139 = _io_exe_rd_0_resp_T_138 | _io_exe_rd_0_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_140 = _io_exe_rd_0_resp_T_139 | _io_exe_rd_0_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_141 = _io_exe_rd_0_resp_T_140 | _io_exe_rd_0_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_142 = _io_exe_rd_0_resp_T_141 | _io_exe_rd_0_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_143 = _io_exe_rd_0_resp_T_142 | _io_exe_rd_0_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_144 = _io_exe_rd_0_resp_T_143 | _io_exe_rd_0_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_145 = _io_exe_rd_0_resp_T_144 | _io_exe_rd_0_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_146 = _io_exe_rd_0_resp_T_145 | _io_exe_rd_0_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_147 = _io_exe_rd_0_resp_T_146 | _io_exe_rd_0_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_148 = _io_exe_rd_0_resp_T_147 | _io_exe_rd_0_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_149 = _io_exe_rd_0_resp_T_148 | _io_exe_rd_0_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_150 = _io_exe_rd_0_resp_T_149 | _io_exe_rd_0_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_0_resp_T_151 = _io_exe_rd_0_resp_T_150 | _io_exe_rd_0_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_1 = io_exe_rd_1_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_8_out_coef_out_1_0 = io_exe_rd_1_req_sel ? io_coef_in_mainch_drc_smooth_2 :
    io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_8_out_coef_out_1_1 = io_exe_rd_1_req_sel ? io_coef_in_mainch_drc_smooth_3 :
    io_coef_in_mainch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_998 = io_exe_rd_1_req_gidx[0] ? tmp_8_out_coef_out_1_1 : tmp_8_out_coef_out_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h2 ? _GEN_998 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_1 = io_exe_rd_1_req_iscoef ? tmp_8_out_out_out_1 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_9_out_coef_out_1_0 = io_exe_rd_1_req_sel ? io_coef_in_subch_drc_smooth_2 :
    io_coef_in_subch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_9_out_coef_out_1_1 = io_exe_rd_1_req_sel ? io_coef_in_subch_drc_smooth_3 :
    io_coef_in_subch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_1002 = io_exe_rd_1_req_gidx[0] ? tmp_9_out_coef_out_1_1 : tmp_9_out_coef_out_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h2 ? _GEN_1002 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_1 = io_exe_rd_1_req_iscoef ? tmp_9_out_out_out_1 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1006 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1007 = 3'h2 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1006; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1008 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1007; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1009 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1008; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1009 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_1 = io_exe_rd_1_req_iscoef ? tmp_10_out_out_out_1 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_1 = io_exe_rd_1_req_iscoef ? tmp_10_out_out_out_1 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1020 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1021 = 3'h2 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1020; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1022 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1021; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1023 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1022; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1023 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_1 = io_exe_rd_1_req_iscoef ? tmp_12_out_out_out_1 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_1 = io_exe_rd_1_req_iscoef ? tmp_12_out_out_out_1 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1034 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1035 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_1034; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1036 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_1035; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1037 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_1036; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1037 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_6 = io_exe_rd_1_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_1040 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1041 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt__2 : _GEN_1040; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1042 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt__3 : _GEN_1041; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1042 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_14_out_out_out_3 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_1 = io_exe_rd_1_req_iscoef ? tmp_14_out_out_out_2 : tmp_14_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1047 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1048 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_1047; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1049 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_1048; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1050 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_1049; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1050 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1053 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1054 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_1_2 : _GEN_1053; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1055 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_1_3 : _GEN_1054; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1055 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_15_out_out_out_3 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_1 = io_exe_rd_1_req_iscoef ? tmp_15_out_out_out_2 : tmp_15_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1060 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1061 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_1060; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1062 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_1061; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1063 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_1062; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1063 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1066 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1067 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_2_2 : _GEN_1066; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1068 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_2_3 : _GEN_1067; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1068 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_16_out_out_out_3 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_1 = io_exe_rd_1_req_iscoef ? tmp_16_out_out_out_2 : tmp_16_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1073 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1074 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_1073; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1075 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_1074; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1076 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_1075; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1076 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1079 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1080 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_3_2 : _GEN_1079; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1081 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_3_3 : _GEN_1080; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1081 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_17_out_out_out_3 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_1 = io_exe_rd_1_req_iscoef ? tmp_17_out_out_out_2 : tmp_17_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1086 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1087 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_1086; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1088 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_1087; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1089 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_1088; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1089 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1092 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1093 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_4_2 : _GEN_1092; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1094 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_4_3 : _GEN_1093; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1094 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_18_out_out_out_3 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_1 = io_exe_rd_1_req_iscoef ? tmp_18_out_out_out_2 : tmp_18_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1099 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1100 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_1099; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1101 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_1100; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1102 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_1101; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1102 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1105 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1106 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_5_2 : _GEN_1105; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1107 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_5_3 : _GEN_1106; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1107 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_19_out_out_out_3 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_1 = io_exe_rd_1_req_iscoef ? tmp_19_out_out_out_2 : tmp_19_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1112 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1113 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_1112; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1114 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_1113; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1115 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_1114; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1115 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1118 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1119 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_6_2 : _GEN_1118; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1120 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_6_3 : _GEN_1119; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1120 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_20_out_out_out_3 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_1 = io_exe_rd_1_req_iscoef ? tmp_20_out_out_out_2 : tmp_20_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1125 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1126 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_1125; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1127 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_1126; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1128 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_1127; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1128 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1131 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1132 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_7_2 : _GEN_1131; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1133 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_7_3 : _GEN_1132; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1133 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_21_out_out_out_3 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_1 = io_exe_rd_1_req_iscoef ? tmp_21_out_out_out_2 : tmp_21_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1138 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1139 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_1138; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1140 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_1139; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1141 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_1140; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1141 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1144 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1145 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_8_2 : _GEN_1144; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1146 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_8_3 : _GEN_1145; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1146 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_22_out_out_out_3 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_1 = io_exe_rd_1_req_iscoef ? tmp_22_out_out_out_2 : tmp_22_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1151 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1152 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_1151; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1153 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_1152; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1154 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_1153; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1154 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1157 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1158 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_9_2 : _GEN_1157; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1159 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_9_3 : _GEN_1158; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1159 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_23_out_out_out_3 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_1 = io_exe_rd_1_req_iscoef ? tmp_23_out_out_out_2 : tmp_23_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1164 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1165 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_1164; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1166 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_1165; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1167 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_1166; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1167 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1170 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1171 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_10_2 : _GEN_1170; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1172 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_10_3 : _GEN_1171; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1172 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_24_out_out_out_3 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_1 = io_exe_rd_1_req_iscoef ? tmp_24_out_out_out_2 : tmp_24_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1177 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1178 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_1177; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1179 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_1178; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1180 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_1179; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1180 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1183 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1184 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_11_2 : _GEN_1183; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1185 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_11_3 : _GEN_1184; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1185 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_25_out_out_out_3 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_1 = io_exe_rd_1_req_iscoef ? tmp_25_out_out_out_2 : tmp_25_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1190 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1191 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_1190; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1192 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_1191; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1193 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_1192; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1193 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1196 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1197 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_12_2 : _GEN_1196; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1198 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_12_3 : _GEN_1197; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1198 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_26_out_out_out_3 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_1 = io_exe_rd_1_req_iscoef ? tmp_26_out_out_out_2 : tmp_26_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1203 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1204 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_1203; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1205 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_1204; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1206 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_1205; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1206 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1209 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1210 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_13_2 : _GEN_1209; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1211 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_13_3 : _GEN_1210; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1211 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_27_out_out_out_3 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_1 = io_exe_rd_1_req_iscoef ? tmp_27_out_out_out_2 : tmp_27_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1216 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1217 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_1216; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1218 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_1217; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1219 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_1218; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1219 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1222 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1223 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_14_2 : _GEN_1222; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1224 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_14_3 : _GEN_1223; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1224 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_28_out_out_out_3 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_1 = io_exe_rd_1_req_iscoef ? tmp_28_out_out_out_2 : tmp_28_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1229 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1230 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_1229; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1231 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_1230; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1232 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_1231; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1232 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1235 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1236 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_15_2 : _GEN_1235; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1237 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_15_3 : _GEN_1236; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1237 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_29_out_out_out_3 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_1 = io_exe_rd_1_req_iscoef ? tmp_29_out_out_out_2 : tmp_29_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1242 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1243 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_1242; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1244 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_1243; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1245 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_1244; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1245 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1248 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1249 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_16_2 : _GEN_1248; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1250 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_16_3 : _GEN_1249; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1250 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_30_out_out_out_3 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_1 = io_exe_rd_1_req_iscoef ? tmp_30_out_out_out_2 : tmp_30_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1255 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1256 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_1255; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1257 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_1256; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1258 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_1257; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1258 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1261 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1262 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_17_2 : _GEN_1261; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1263 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_17_3 : _GEN_1262; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1263 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_31_out_out_out_3 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_1 = io_exe_rd_1_req_iscoef ? tmp_31_out_out_out_2 : tmp_31_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1268 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1269 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_1268; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1270 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_1269; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1271 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_1270; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1271 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1274 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1275 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_18_2 : _GEN_1274; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1276 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_18_3 : _GEN_1275; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1276 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_32_out_out_out_3 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_1 = io_exe_rd_1_req_iscoef ? tmp_32_out_out_out_2 : tmp_32_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1281 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1282 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_1281; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1283 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_1282; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1284 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_1283; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1284 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1287 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1288 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_19_2 : _GEN_1287; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1289 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_19_3 : _GEN_1288; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1289 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_33_out_out_out_3 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_1 = io_exe_rd_1_req_iscoef ? tmp_33_out_out_out_2 : tmp_33_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1294 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1295 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_1294; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1296 = 3'h3 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_1295; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1297 = 3'h4 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_1296; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_2 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1297 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1300 = 2'h1 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1301 = 2'h2 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_20_2 : _GEN_1300; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1302 = 2'h3 == _tmp_14_out_out_T_6[1:0] ? reg_type5_data_nxt_20_3 : _GEN_1301; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_3 = _tmp_14_out_out_T_6 < 3'h4 ? _GEN_1302 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_3 = io_exe_rd_1_req_isgroup ? tmp_34_out_out_out_3 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_1 = io_exe_rd_1_req_iscoef ? tmp_34_out_out_out_2 : tmp_34_out_out_3; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1307 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1308 = 3'h2 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1307; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1309 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1308; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1310 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1309; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1310 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_1 = io_exe_rd_1_req_iscoef ? tmp_35_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1314 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1315 = 3'h2 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1314; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1316 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1315; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1317 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1316; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1317 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_1 = io_exe_rd_1_req_iscoef ? tmp_36_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1321 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1322 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_1321; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1323 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1322; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1324 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1323; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1324 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_1 = io_exe_rd_1_req_iscoef ? tmp_37_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1328 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1329 = 3'h2 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1328; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1330 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1329; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1331 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1330; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1331 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_1 = io_exe_rd_1_req_iscoef ? tmp_38_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1335 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1336 = 3'h2 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1335; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1337 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1336; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1338 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1337; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1338 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_1 = io_exe_rd_1_req_iscoef ? tmp_39_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1342 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1343 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_1342; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1344 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1343; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1345 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1344; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1345 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_1 = io_exe_rd_1_req_iscoef ? tmp_40_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1349 = 3'h1 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1350 = 3'h2 == io_exe_rd_1_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_1349; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1351 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1350; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1352 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1351; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1352 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_1 = io_exe_rd_1_req_iscoef ? tmp_41_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1356 = 3'h1 == io_exe_rd_1_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1357 = 3'h2 == io_exe_rd_1_req_gidx ? reg_type6_coef_7_2 : _GEN_1356; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1358 = 3'h3 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1357; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1359 = 3'h4 == io_exe_rd_1_req_gidx ? 32'h0 : _GEN_1358; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_1 = io_exe_rd_1_req_gidx < 3'h5 ? _GEN_1359 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_1 = io_exe_rd_1_req_iscoef ? tmp_42_out_out_out_1 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_1 = io_exe_rd_1_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_1 = io_exe_rd_1_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_1 = io_exe_rd_1_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_1 = io_exe_rd_1_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_1 = io_exe_rd_1_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_1 = io_exe_rd_1_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_1 = io_exe_rd_1_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_1 = io_exe_rd_1_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_1_resp_T = 64'h1 << io_exe_rd_1_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_1_resp_T_52 = _io_exe_rd_1_resp_T[0] ? tmp_0_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_53 = _io_exe_rd_1_resp_T[1] ? tmp_1_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_54 = _io_exe_rd_1_resp_T[2] ? tmp_2_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_55 = _io_exe_rd_1_resp_T[3] ? tmp_3_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_56 = _io_exe_rd_1_resp_T[4] ? tmp_4_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_57 = _io_exe_rd_1_resp_T[5] ? tmp_5_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_58 = _io_exe_rd_1_resp_T[6] ? tmp_6_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_59 = _io_exe_rd_1_resp_T[7] ? tmp_7_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_60 = _io_exe_rd_1_resp_T[8] ? tmp_8_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_61 = _io_exe_rd_1_resp_T[9] ? tmp_9_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_62 = _io_exe_rd_1_resp_T[10] ? tmp_10_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_63 = _io_exe_rd_1_resp_T[11] ? tmp_11_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_64 = _io_exe_rd_1_resp_T[12] ? tmp_12_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_65 = _io_exe_rd_1_resp_T[13] ? tmp_13_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_66 = _io_exe_rd_1_resp_T[14] ? tmp_14_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_67 = _io_exe_rd_1_resp_T[15] ? tmp_15_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_68 = _io_exe_rd_1_resp_T[16] ? tmp_16_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_69 = _io_exe_rd_1_resp_T[17] ? tmp_17_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_70 = _io_exe_rd_1_resp_T[18] ? tmp_18_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_71 = _io_exe_rd_1_resp_T[19] ? tmp_19_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_72 = _io_exe_rd_1_resp_T[20] ? tmp_20_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_73 = _io_exe_rd_1_resp_T[21] ? tmp_21_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_74 = _io_exe_rd_1_resp_T[22] ? tmp_22_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_75 = _io_exe_rd_1_resp_T[23] ? tmp_23_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_76 = _io_exe_rd_1_resp_T[24] ? tmp_24_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_77 = _io_exe_rd_1_resp_T[25] ? tmp_25_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_78 = _io_exe_rd_1_resp_T[26] ? tmp_26_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_79 = _io_exe_rd_1_resp_T[27] ? tmp_27_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_80 = _io_exe_rd_1_resp_T[28] ? tmp_28_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_81 = _io_exe_rd_1_resp_T[29] ? tmp_29_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_82 = _io_exe_rd_1_resp_T[30] ? tmp_30_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_83 = _io_exe_rd_1_resp_T[31] ? tmp_31_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_84 = _io_exe_rd_1_resp_T[32] ? tmp_32_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_85 = _io_exe_rd_1_resp_T[33] ? tmp_33_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_86 = _io_exe_rd_1_resp_T[34] ? tmp_34_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_87 = _io_exe_rd_1_resp_T[35] ? tmp_35_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_88 = _io_exe_rd_1_resp_T[36] ? tmp_36_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_89 = _io_exe_rd_1_resp_T[37] ? tmp_37_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_90 = _io_exe_rd_1_resp_T[38] ? tmp_38_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_91 = _io_exe_rd_1_resp_T[39] ? tmp_39_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_92 = _io_exe_rd_1_resp_T[40] ? tmp_40_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_93 = _io_exe_rd_1_resp_T[41] ? tmp_41_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_94 = _io_exe_rd_1_resp_T[42] ? tmp_42_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_95 = _io_exe_rd_1_resp_T[43] ? tmp_43_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_96 = _io_exe_rd_1_resp_T[44] ? tmp_44_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_97 = _io_exe_rd_1_resp_T[45] ? tmp_45_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_98 = _io_exe_rd_1_resp_T[46] ? tmp_46_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_99 = _io_exe_rd_1_resp_T[47] ? tmp_47_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_100 = _io_exe_rd_1_resp_T[48] ? tmp_48_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_101 = _io_exe_rd_1_resp_T[49] ? tmp_49_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_102 = _io_exe_rd_1_resp_T[50] ? tmp_50_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_103 = _io_exe_rd_1_resp_T_52 | _io_exe_rd_1_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_104 = _io_exe_rd_1_resp_T_103 | _io_exe_rd_1_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_105 = _io_exe_rd_1_resp_T_104 | _io_exe_rd_1_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_106 = _io_exe_rd_1_resp_T_105 | _io_exe_rd_1_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_107 = _io_exe_rd_1_resp_T_106 | _io_exe_rd_1_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_108 = _io_exe_rd_1_resp_T_107 | _io_exe_rd_1_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_109 = _io_exe_rd_1_resp_T_108 | _io_exe_rd_1_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_110 = _io_exe_rd_1_resp_T_109 | _io_exe_rd_1_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_111 = _io_exe_rd_1_resp_T_110 | _io_exe_rd_1_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_112 = _io_exe_rd_1_resp_T_111 | _io_exe_rd_1_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_113 = _io_exe_rd_1_resp_T_112 | _io_exe_rd_1_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_114 = _io_exe_rd_1_resp_T_113 | _io_exe_rd_1_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_115 = _io_exe_rd_1_resp_T_114 | _io_exe_rd_1_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_116 = _io_exe_rd_1_resp_T_115 | _io_exe_rd_1_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_117 = _io_exe_rd_1_resp_T_116 | _io_exe_rd_1_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_118 = _io_exe_rd_1_resp_T_117 | _io_exe_rd_1_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_119 = _io_exe_rd_1_resp_T_118 | _io_exe_rd_1_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_120 = _io_exe_rd_1_resp_T_119 | _io_exe_rd_1_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_121 = _io_exe_rd_1_resp_T_120 | _io_exe_rd_1_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_122 = _io_exe_rd_1_resp_T_121 | _io_exe_rd_1_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_123 = _io_exe_rd_1_resp_T_122 | _io_exe_rd_1_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_124 = _io_exe_rd_1_resp_T_123 | _io_exe_rd_1_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_125 = _io_exe_rd_1_resp_T_124 | _io_exe_rd_1_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_126 = _io_exe_rd_1_resp_T_125 | _io_exe_rd_1_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_127 = _io_exe_rd_1_resp_T_126 | _io_exe_rd_1_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_128 = _io_exe_rd_1_resp_T_127 | _io_exe_rd_1_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_129 = _io_exe_rd_1_resp_T_128 | _io_exe_rd_1_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_130 = _io_exe_rd_1_resp_T_129 | _io_exe_rd_1_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_131 = _io_exe_rd_1_resp_T_130 | _io_exe_rd_1_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_132 = _io_exe_rd_1_resp_T_131 | _io_exe_rd_1_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_133 = _io_exe_rd_1_resp_T_132 | _io_exe_rd_1_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_134 = _io_exe_rd_1_resp_T_133 | _io_exe_rd_1_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_135 = _io_exe_rd_1_resp_T_134 | _io_exe_rd_1_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_136 = _io_exe_rd_1_resp_T_135 | _io_exe_rd_1_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_137 = _io_exe_rd_1_resp_T_136 | _io_exe_rd_1_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_138 = _io_exe_rd_1_resp_T_137 | _io_exe_rd_1_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_139 = _io_exe_rd_1_resp_T_138 | _io_exe_rd_1_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_140 = _io_exe_rd_1_resp_T_139 | _io_exe_rd_1_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_141 = _io_exe_rd_1_resp_T_140 | _io_exe_rd_1_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_142 = _io_exe_rd_1_resp_T_141 | _io_exe_rd_1_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_143 = _io_exe_rd_1_resp_T_142 | _io_exe_rd_1_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_144 = _io_exe_rd_1_resp_T_143 | _io_exe_rd_1_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_145 = _io_exe_rd_1_resp_T_144 | _io_exe_rd_1_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_146 = _io_exe_rd_1_resp_T_145 | _io_exe_rd_1_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_147 = _io_exe_rd_1_resp_T_146 | _io_exe_rd_1_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_148 = _io_exe_rd_1_resp_T_147 | _io_exe_rd_1_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_149 = _io_exe_rd_1_resp_T_148 | _io_exe_rd_1_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_150 = _io_exe_rd_1_resp_T_149 | _io_exe_rd_1_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_1_resp_T_151 = _io_exe_rd_1_resp_T_150 | _io_exe_rd_1_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_2 = io_exe_rd_2_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1379 = io_exe_rd_2_req_gidx[0] ? io_coef_in_mainch_drc_smooth_1 : io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h2 ? _GEN_1379 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_2 = io_exe_rd_2_req_iscoef ? tmp_8_out_out_out_2 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1383 = io_exe_rd_2_req_gidx[0] ? io_coef_in_subch_drc_smooth_1 : io_coef_in_subch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h2 ? _GEN_1383 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_2 = io_exe_rd_2_req_iscoef ? tmp_9_out_out_out_2 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1387 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1388 = 3'h2 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1387; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1389 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1388; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1390 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1389; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1390 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_2 = io_exe_rd_2_req_iscoef ? tmp_10_out_out_out_2 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_2 = io_exe_rd_2_req_iscoef ? tmp_10_out_out_out_2 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1401 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1402 = 3'h2 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1401; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1403 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1402; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1404 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1403; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1404 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_2 = io_exe_rd_2_req_iscoef ? tmp_12_out_out_out_2 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_2 = io_exe_rd_2_req_iscoef ? tmp_12_out_out_out_2 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1415 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1416 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_1415; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1417 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_1416; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1418 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_1417; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1418 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_10 = io_exe_rd_2_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_1421 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1422 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt__2 : _GEN_1421; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1423 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt__3 : _GEN_1422; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1423 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_14_out_out_out_5 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_2 = io_exe_rd_2_req_iscoef ? tmp_14_out_out_out_4 : tmp_14_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1428 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1429 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_1428; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1430 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_1429; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1431 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_1430; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1431 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1434 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1435 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_1_2 : _GEN_1434; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1436 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_1_3 : _GEN_1435; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1436 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_15_out_out_out_5 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_2 = io_exe_rd_2_req_iscoef ? tmp_15_out_out_out_4 : tmp_15_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1441 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1442 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_1441; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1443 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_1442; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1444 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_1443; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1444 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1447 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1448 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_2_2 : _GEN_1447; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1449 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_2_3 : _GEN_1448; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1449 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_16_out_out_out_5 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_2 = io_exe_rd_2_req_iscoef ? tmp_16_out_out_out_4 : tmp_16_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1454 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1455 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_1454; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1456 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_1455; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1457 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_1456; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1457 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1460 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1461 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_3_2 : _GEN_1460; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1462 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_3_3 : _GEN_1461; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1462 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_17_out_out_out_5 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_2 = io_exe_rd_2_req_iscoef ? tmp_17_out_out_out_4 : tmp_17_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1467 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1468 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_1467; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1469 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_1468; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1470 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_1469; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1470 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1473 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1474 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_4_2 : _GEN_1473; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1475 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_4_3 : _GEN_1474; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1475 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_18_out_out_out_5 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_2 = io_exe_rd_2_req_iscoef ? tmp_18_out_out_out_4 : tmp_18_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1480 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1481 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_1480; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1482 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_1481; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1483 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_1482; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1483 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1486 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1487 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_5_2 : _GEN_1486; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1488 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_5_3 : _GEN_1487; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1488 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_19_out_out_out_5 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_2 = io_exe_rd_2_req_iscoef ? tmp_19_out_out_out_4 : tmp_19_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1493 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1494 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_1493; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1495 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_1494; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1496 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_1495; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1496 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1499 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1500 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_6_2 : _GEN_1499; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1501 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_6_3 : _GEN_1500; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1501 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_20_out_out_out_5 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_2 = io_exe_rd_2_req_iscoef ? tmp_20_out_out_out_4 : tmp_20_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1506 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1507 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_1506; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1508 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_1507; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1509 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_1508; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1509 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1512 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1513 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_7_2 : _GEN_1512; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1514 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_7_3 : _GEN_1513; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1514 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_21_out_out_out_5 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_2 = io_exe_rd_2_req_iscoef ? tmp_21_out_out_out_4 : tmp_21_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1519 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1520 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_1519; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1521 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_1520; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1522 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_1521; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1522 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1525 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1526 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_8_2 : _GEN_1525; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1527 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_8_3 : _GEN_1526; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1527 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_22_out_out_out_5 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_2 = io_exe_rd_2_req_iscoef ? tmp_22_out_out_out_4 : tmp_22_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1532 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1533 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_1532; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1534 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_1533; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1535 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_1534; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1535 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1538 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1539 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_9_2 : _GEN_1538; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1540 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_9_3 : _GEN_1539; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1540 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_23_out_out_out_5 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_2 = io_exe_rd_2_req_iscoef ? tmp_23_out_out_out_4 : tmp_23_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1545 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1546 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_1545; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1547 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_1546; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1548 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_1547; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1548 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1551 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1552 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_10_2 : _GEN_1551; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1553 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_10_3 : _GEN_1552; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1553 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_24_out_out_out_5 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_2 = io_exe_rd_2_req_iscoef ? tmp_24_out_out_out_4 : tmp_24_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1558 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1559 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_1558; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1560 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_1559; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1561 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_1560; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1561 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1564 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1565 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_11_2 : _GEN_1564; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1566 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_11_3 : _GEN_1565; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1566 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_25_out_out_out_5 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_2 = io_exe_rd_2_req_iscoef ? tmp_25_out_out_out_4 : tmp_25_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1571 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1572 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_1571; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1573 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_1572; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1574 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_1573; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1574 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1577 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1578 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_12_2 : _GEN_1577; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1579 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_12_3 : _GEN_1578; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1579 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_26_out_out_out_5 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_2 = io_exe_rd_2_req_iscoef ? tmp_26_out_out_out_4 : tmp_26_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1584 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1585 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_1584; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1586 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_1585; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1587 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_1586; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1587 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1590 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1591 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_13_2 : _GEN_1590; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1592 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_13_3 : _GEN_1591; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1592 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_27_out_out_out_5 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_2 = io_exe_rd_2_req_iscoef ? tmp_27_out_out_out_4 : tmp_27_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1597 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1598 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_1597; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1599 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_1598; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1600 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_1599; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1600 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1603 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1604 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_14_2 : _GEN_1603; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1605 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_14_3 : _GEN_1604; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1605 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_28_out_out_out_5 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_2 = io_exe_rd_2_req_iscoef ? tmp_28_out_out_out_4 : tmp_28_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1610 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1611 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_1610; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1612 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_1611; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1613 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_1612; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1613 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1616 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1617 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_15_2 : _GEN_1616; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1618 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_15_3 : _GEN_1617; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1618 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_29_out_out_out_5 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_2 = io_exe_rd_2_req_iscoef ? tmp_29_out_out_out_4 : tmp_29_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1623 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1624 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_1623; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1625 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_1624; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1626 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_1625; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1626 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1629 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1630 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_16_2 : _GEN_1629; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1631 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_16_3 : _GEN_1630; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1631 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_30_out_out_out_5 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_2 = io_exe_rd_2_req_iscoef ? tmp_30_out_out_out_4 : tmp_30_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1636 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1637 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_1636; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1638 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_1637; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1639 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_1638; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1639 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1642 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1643 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_17_2 : _GEN_1642; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1644 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_17_3 : _GEN_1643; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1644 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_31_out_out_out_5 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_2 = io_exe_rd_2_req_iscoef ? tmp_31_out_out_out_4 : tmp_31_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1649 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1650 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_1649; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1651 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_1650; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1652 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_1651; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1652 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1655 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1656 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_18_2 : _GEN_1655; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1657 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_18_3 : _GEN_1656; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1657 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_32_out_out_out_5 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_2 = io_exe_rd_2_req_iscoef ? tmp_32_out_out_out_4 : tmp_32_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1662 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1663 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_1662; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1664 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_1663; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1665 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_1664; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1665 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1668 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1669 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_19_2 : _GEN_1668; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1670 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_19_3 : _GEN_1669; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1670 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_33_out_out_out_5 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_2 = io_exe_rd_2_req_iscoef ? tmp_33_out_out_out_4 : tmp_33_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1675 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1676 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_1675; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1677 = 3'h3 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_1676; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1678 = 3'h4 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_1677; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_4 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1678 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1681 = 2'h1 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1682 = 2'h2 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_20_2 : _GEN_1681; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1683 = 2'h3 == _tmp_14_out_out_T_10[1:0] ? reg_type5_data_nxt_20_3 : _GEN_1682; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_5 = _tmp_14_out_out_T_10 < 3'h4 ? _GEN_1683 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_5 = io_exe_rd_2_req_isgroup ? tmp_34_out_out_out_5 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_2 = io_exe_rd_2_req_iscoef ? tmp_34_out_out_out_4 : tmp_34_out_out_5; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1688 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1689 = 3'h2 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1688; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1690 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1689; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1691 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1690; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1691 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_2 = io_exe_rd_2_req_iscoef ? tmp_35_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1695 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1696 = 3'h2 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1695; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1697 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1696; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1698 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1697; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1698 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_2 = io_exe_rd_2_req_iscoef ? tmp_36_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1702 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1703 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_1702; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1704 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1703; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1705 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1704; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1705 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_2 = io_exe_rd_2_req_iscoef ? tmp_37_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1709 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1710 = 3'h2 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1709; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1711 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1710; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1712 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1711; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1712 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_2 = io_exe_rd_2_req_iscoef ? tmp_38_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1716 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1717 = 3'h2 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1716; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1718 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1717; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1719 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1718; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1719 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_2 = io_exe_rd_2_req_iscoef ? tmp_39_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1723 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1724 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_1723; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1725 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1724; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1726 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1725; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1726 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_2 = io_exe_rd_2_req_iscoef ? tmp_40_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1730 = 3'h1 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1731 = 3'h2 == io_exe_rd_2_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_1730; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1732 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1731; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1733 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1732; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1733 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_2 = io_exe_rd_2_req_iscoef ? tmp_41_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1737 = 3'h1 == io_exe_rd_2_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1738 = 3'h2 == io_exe_rd_2_req_gidx ? reg_type6_coef_7_2 : _GEN_1737; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1739 = 3'h3 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1738; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1740 = 3'h4 == io_exe_rd_2_req_gidx ? 32'h0 : _GEN_1739; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_2 = io_exe_rd_2_req_gidx < 3'h5 ? _GEN_1740 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_2 = io_exe_rd_2_req_iscoef ? tmp_42_out_out_out_2 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_2 = io_exe_rd_2_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_2 = io_exe_rd_2_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_2 = io_exe_rd_2_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_2 = io_exe_rd_2_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_2 = io_exe_rd_2_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_2 = io_exe_rd_2_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_2 = io_exe_rd_2_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_2 = io_exe_rd_2_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_2_resp_T = 64'h1 << io_exe_rd_2_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_2_resp_T_52 = _io_exe_rd_2_resp_T[0] ? tmp_0_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_53 = _io_exe_rd_2_resp_T[1] ? tmp_1_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_54 = _io_exe_rd_2_resp_T[2] ? tmp_2_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_55 = _io_exe_rd_2_resp_T[3] ? tmp_3_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_56 = _io_exe_rd_2_resp_T[4] ? tmp_4_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_57 = _io_exe_rd_2_resp_T[5] ? tmp_5_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_58 = _io_exe_rd_2_resp_T[6] ? tmp_6_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_59 = _io_exe_rd_2_resp_T[7] ? tmp_7_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_60 = _io_exe_rd_2_resp_T[8] ? tmp_8_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_61 = _io_exe_rd_2_resp_T[9] ? tmp_9_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_62 = _io_exe_rd_2_resp_T[10] ? tmp_10_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_63 = _io_exe_rd_2_resp_T[11] ? tmp_11_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_64 = _io_exe_rd_2_resp_T[12] ? tmp_12_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_65 = _io_exe_rd_2_resp_T[13] ? tmp_13_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_66 = _io_exe_rd_2_resp_T[14] ? tmp_14_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_67 = _io_exe_rd_2_resp_T[15] ? tmp_15_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_68 = _io_exe_rd_2_resp_T[16] ? tmp_16_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_69 = _io_exe_rd_2_resp_T[17] ? tmp_17_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_70 = _io_exe_rd_2_resp_T[18] ? tmp_18_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_71 = _io_exe_rd_2_resp_T[19] ? tmp_19_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_72 = _io_exe_rd_2_resp_T[20] ? tmp_20_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_73 = _io_exe_rd_2_resp_T[21] ? tmp_21_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_74 = _io_exe_rd_2_resp_T[22] ? tmp_22_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_75 = _io_exe_rd_2_resp_T[23] ? tmp_23_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_76 = _io_exe_rd_2_resp_T[24] ? tmp_24_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_77 = _io_exe_rd_2_resp_T[25] ? tmp_25_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_78 = _io_exe_rd_2_resp_T[26] ? tmp_26_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_79 = _io_exe_rd_2_resp_T[27] ? tmp_27_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_80 = _io_exe_rd_2_resp_T[28] ? tmp_28_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_81 = _io_exe_rd_2_resp_T[29] ? tmp_29_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_82 = _io_exe_rd_2_resp_T[30] ? tmp_30_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_83 = _io_exe_rd_2_resp_T[31] ? tmp_31_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_84 = _io_exe_rd_2_resp_T[32] ? tmp_32_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_85 = _io_exe_rd_2_resp_T[33] ? tmp_33_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_86 = _io_exe_rd_2_resp_T[34] ? tmp_34_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_87 = _io_exe_rd_2_resp_T[35] ? tmp_35_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_88 = _io_exe_rd_2_resp_T[36] ? tmp_36_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_89 = _io_exe_rd_2_resp_T[37] ? tmp_37_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_90 = _io_exe_rd_2_resp_T[38] ? tmp_38_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_91 = _io_exe_rd_2_resp_T[39] ? tmp_39_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_92 = _io_exe_rd_2_resp_T[40] ? tmp_40_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_93 = _io_exe_rd_2_resp_T[41] ? tmp_41_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_94 = _io_exe_rd_2_resp_T[42] ? tmp_42_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_95 = _io_exe_rd_2_resp_T[43] ? tmp_43_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_96 = _io_exe_rd_2_resp_T[44] ? tmp_44_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_97 = _io_exe_rd_2_resp_T[45] ? tmp_45_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_98 = _io_exe_rd_2_resp_T[46] ? tmp_46_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_99 = _io_exe_rd_2_resp_T[47] ? tmp_47_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_100 = _io_exe_rd_2_resp_T[48] ? tmp_48_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_101 = _io_exe_rd_2_resp_T[49] ? tmp_49_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_102 = _io_exe_rd_2_resp_T[50] ? tmp_50_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_103 = _io_exe_rd_2_resp_T_52 | _io_exe_rd_2_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_104 = _io_exe_rd_2_resp_T_103 | _io_exe_rd_2_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_105 = _io_exe_rd_2_resp_T_104 | _io_exe_rd_2_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_106 = _io_exe_rd_2_resp_T_105 | _io_exe_rd_2_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_107 = _io_exe_rd_2_resp_T_106 | _io_exe_rd_2_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_108 = _io_exe_rd_2_resp_T_107 | _io_exe_rd_2_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_109 = _io_exe_rd_2_resp_T_108 | _io_exe_rd_2_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_110 = _io_exe_rd_2_resp_T_109 | _io_exe_rd_2_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_111 = _io_exe_rd_2_resp_T_110 | _io_exe_rd_2_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_112 = _io_exe_rd_2_resp_T_111 | _io_exe_rd_2_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_113 = _io_exe_rd_2_resp_T_112 | _io_exe_rd_2_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_114 = _io_exe_rd_2_resp_T_113 | _io_exe_rd_2_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_115 = _io_exe_rd_2_resp_T_114 | _io_exe_rd_2_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_116 = _io_exe_rd_2_resp_T_115 | _io_exe_rd_2_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_117 = _io_exe_rd_2_resp_T_116 | _io_exe_rd_2_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_118 = _io_exe_rd_2_resp_T_117 | _io_exe_rd_2_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_119 = _io_exe_rd_2_resp_T_118 | _io_exe_rd_2_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_120 = _io_exe_rd_2_resp_T_119 | _io_exe_rd_2_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_121 = _io_exe_rd_2_resp_T_120 | _io_exe_rd_2_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_122 = _io_exe_rd_2_resp_T_121 | _io_exe_rd_2_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_123 = _io_exe_rd_2_resp_T_122 | _io_exe_rd_2_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_124 = _io_exe_rd_2_resp_T_123 | _io_exe_rd_2_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_125 = _io_exe_rd_2_resp_T_124 | _io_exe_rd_2_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_126 = _io_exe_rd_2_resp_T_125 | _io_exe_rd_2_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_127 = _io_exe_rd_2_resp_T_126 | _io_exe_rd_2_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_128 = _io_exe_rd_2_resp_T_127 | _io_exe_rd_2_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_129 = _io_exe_rd_2_resp_T_128 | _io_exe_rd_2_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_130 = _io_exe_rd_2_resp_T_129 | _io_exe_rd_2_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_131 = _io_exe_rd_2_resp_T_130 | _io_exe_rd_2_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_132 = _io_exe_rd_2_resp_T_131 | _io_exe_rd_2_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_133 = _io_exe_rd_2_resp_T_132 | _io_exe_rd_2_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_134 = _io_exe_rd_2_resp_T_133 | _io_exe_rd_2_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_135 = _io_exe_rd_2_resp_T_134 | _io_exe_rd_2_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_136 = _io_exe_rd_2_resp_T_135 | _io_exe_rd_2_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_137 = _io_exe_rd_2_resp_T_136 | _io_exe_rd_2_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_138 = _io_exe_rd_2_resp_T_137 | _io_exe_rd_2_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_139 = _io_exe_rd_2_resp_T_138 | _io_exe_rd_2_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_140 = _io_exe_rd_2_resp_T_139 | _io_exe_rd_2_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_141 = _io_exe_rd_2_resp_T_140 | _io_exe_rd_2_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_142 = _io_exe_rd_2_resp_T_141 | _io_exe_rd_2_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_143 = _io_exe_rd_2_resp_T_142 | _io_exe_rd_2_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_144 = _io_exe_rd_2_resp_T_143 | _io_exe_rd_2_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_145 = _io_exe_rd_2_resp_T_144 | _io_exe_rd_2_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_146 = _io_exe_rd_2_resp_T_145 | _io_exe_rd_2_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_147 = _io_exe_rd_2_resp_T_146 | _io_exe_rd_2_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_148 = _io_exe_rd_2_resp_T_147 | _io_exe_rd_2_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_149 = _io_exe_rd_2_resp_T_148 | _io_exe_rd_2_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_150 = _io_exe_rd_2_resp_T_149 | _io_exe_rd_2_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_2_resp_T_151 = _io_exe_rd_2_resp_T_150 | _io_exe_rd_2_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_3 = io_exe_rd_3_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_8_out_coef_out_3_0 = io_exe_rd_3_req_sel ? io_coef_in_mainch_drc_smooth_2 :
    io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_8_out_coef_out_3_1 = io_exe_rd_3_req_sel ? io_coef_in_mainch_drc_smooth_3 :
    io_coef_in_mainch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_1760 = io_exe_rd_3_req_gidx[0] ? tmp_8_out_coef_out_3_1 : tmp_8_out_coef_out_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h2 ? _GEN_1760 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_3 = io_exe_rd_3_req_iscoef ? tmp_8_out_out_out_3 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_9_out_coef_out_3_0 = io_exe_rd_3_req_sel ? io_coef_in_subch_drc_smooth_2 :
    io_coef_in_subch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_9_out_coef_out_3_1 = io_exe_rd_3_req_sel ? io_coef_in_subch_drc_smooth_3 :
    io_coef_in_subch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_1764 = io_exe_rd_3_req_gidx[0] ? tmp_9_out_coef_out_3_1 : tmp_9_out_coef_out_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h2 ? _GEN_1764 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_3 = io_exe_rd_3_req_iscoef ? tmp_9_out_out_out_3 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1768 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1769 = 3'h2 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_1768; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1770 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_1769; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1771 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_1770; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1771 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_3 = io_exe_rd_3_req_iscoef ? tmp_10_out_out_out_3 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_3 = io_exe_rd_3_req_iscoef ? tmp_10_out_out_out_3 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1782 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1783 = 3'h2 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_1782; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1784 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_1783; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1785 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_1784; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1785 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_3 = io_exe_rd_3_req_iscoef ? tmp_12_out_out_out_3 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_3 = io_exe_rd_3_req_iscoef ? tmp_12_out_out_out_3 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1796 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1797 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_1796; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1798 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_1797; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1799 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_1798; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1799 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_14 = io_exe_rd_3_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_1802 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1803 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt__2 : _GEN_1802; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1804 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt__3 : _GEN_1803; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1804 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_14_out_out_out_7 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_3 = io_exe_rd_3_req_iscoef ? tmp_14_out_out_out_6 : tmp_14_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1809 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1810 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_1809; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1811 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_1810; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1812 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_1811; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1812 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1815 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1816 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_1_2 : _GEN_1815; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1817 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_1_3 : _GEN_1816; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1817 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_15_out_out_out_7 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_3 = io_exe_rd_3_req_iscoef ? tmp_15_out_out_out_6 : tmp_15_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1822 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1823 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_1822; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1824 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_1823; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1825 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_1824; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1825 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1828 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1829 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_2_2 : _GEN_1828; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1830 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_2_3 : _GEN_1829; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1830 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_16_out_out_out_7 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_3 = io_exe_rd_3_req_iscoef ? tmp_16_out_out_out_6 : tmp_16_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1835 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1836 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_1835; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1837 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_1836; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1838 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_1837; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1838 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1841 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1842 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_3_2 : _GEN_1841; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1843 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_3_3 : _GEN_1842; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1843 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_17_out_out_out_7 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_3 = io_exe_rd_3_req_iscoef ? tmp_17_out_out_out_6 : tmp_17_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1848 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1849 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_1848; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1850 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_1849; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1851 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_1850; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1851 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1854 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1855 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_4_2 : _GEN_1854; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1856 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_4_3 : _GEN_1855; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1856 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_18_out_out_out_7 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_3 = io_exe_rd_3_req_iscoef ? tmp_18_out_out_out_6 : tmp_18_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1861 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1862 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_1861; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1863 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_1862; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1864 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_1863; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1864 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1867 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1868 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_5_2 : _GEN_1867; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1869 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_5_3 : _GEN_1868; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1869 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_19_out_out_out_7 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_3 = io_exe_rd_3_req_iscoef ? tmp_19_out_out_out_6 : tmp_19_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1874 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1875 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_1874; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1876 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_1875; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1877 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_1876; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1877 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1880 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1881 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_6_2 : _GEN_1880; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1882 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_6_3 : _GEN_1881; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1882 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_20_out_out_out_7 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_3 = io_exe_rd_3_req_iscoef ? tmp_20_out_out_out_6 : tmp_20_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1887 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1888 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_1887; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1889 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_1888; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1890 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_1889; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1890 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1893 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1894 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_7_2 : _GEN_1893; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1895 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_7_3 : _GEN_1894; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1895 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_21_out_out_out_7 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_3 = io_exe_rd_3_req_iscoef ? tmp_21_out_out_out_6 : tmp_21_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1900 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1901 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_1900; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1902 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_1901; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1903 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_1902; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1903 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1906 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1907 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_8_2 : _GEN_1906; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1908 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_8_3 : _GEN_1907; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1908 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_22_out_out_out_7 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_3 = io_exe_rd_3_req_iscoef ? tmp_22_out_out_out_6 : tmp_22_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1913 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1914 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_1913; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1915 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_1914; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1916 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_1915; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1916 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1919 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1920 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_9_2 : _GEN_1919; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1921 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_9_3 : _GEN_1920; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1921 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_23_out_out_out_7 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_3 = io_exe_rd_3_req_iscoef ? tmp_23_out_out_out_6 : tmp_23_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1926 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1927 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_1926; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1928 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_1927; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1929 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_1928; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1929 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1932 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1933 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_10_2 : _GEN_1932; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1934 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_10_3 : _GEN_1933; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1934 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_24_out_out_out_7 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_3 = io_exe_rd_3_req_iscoef ? tmp_24_out_out_out_6 : tmp_24_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1939 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1940 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_1939; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1941 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_1940; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1942 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_1941; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1942 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1945 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1946 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_11_2 : _GEN_1945; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1947 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_11_3 : _GEN_1946; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1947 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_25_out_out_out_7 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_3 = io_exe_rd_3_req_iscoef ? tmp_25_out_out_out_6 : tmp_25_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1952 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1953 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_1952; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1954 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_1953; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1955 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_1954; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1955 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1958 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1959 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_12_2 : _GEN_1958; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1960 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_12_3 : _GEN_1959; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1960 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_26_out_out_out_7 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_3 = io_exe_rd_3_req_iscoef ? tmp_26_out_out_out_6 : tmp_26_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1965 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1966 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_1965; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1967 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_1966; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1968 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_1967; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1968 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1971 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1972 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_13_2 : _GEN_1971; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1973 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_13_3 : _GEN_1972; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1973 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_27_out_out_out_7 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_3 = io_exe_rd_3_req_iscoef ? tmp_27_out_out_out_6 : tmp_27_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1978 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1979 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_1978; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1980 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_1979; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1981 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_1980; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1981 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1984 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1985 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_14_2 : _GEN_1984; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1986 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_14_3 : _GEN_1985; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1986 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_28_out_out_out_7 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_3 = io_exe_rd_3_req_iscoef ? tmp_28_out_out_out_6 : tmp_28_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_1991 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1992 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_1991; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1993 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_1992; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1994 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_1993; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_1994 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_1997 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1998 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_15_2 : _GEN_1997; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_1999 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_15_3 : _GEN_1998; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_1999 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_29_out_out_out_7 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_3 = io_exe_rd_3_req_iscoef ? tmp_29_out_out_out_6 : tmp_29_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2004 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2005 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_2004; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2006 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_2005; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2007 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_2006; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2007 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2010 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2011 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_16_2 : _GEN_2010; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2012 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_16_3 : _GEN_2011; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_2012 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_30_out_out_out_7 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_3 = io_exe_rd_3_req_iscoef ? tmp_30_out_out_out_6 : tmp_30_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2017 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2018 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_2017; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2019 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_2018; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2020 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_2019; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2020 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2023 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2024 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_17_2 : _GEN_2023; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2025 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_17_3 : _GEN_2024; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_2025 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_31_out_out_out_7 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_3 = io_exe_rd_3_req_iscoef ? tmp_31_out_out_out_6 : tmp_31_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2030 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2031 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_2030; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2032 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_2031; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2033 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_2032; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2033 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2036 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2037 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_18_2 : _GEN_2036; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2038 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_18_3 : _GEN_2037; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_2038 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_32_out_out_out_7 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_3 = io_exe_rd_3_req_iscoef ? tmp_32_out_out_out_6 : tmp_32_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2043 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2044 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_2043; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2045 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_2044; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2046 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_2045; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2046 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2049 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2050 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_19_2 : _GEN_2049; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2051 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_19_3 : _GEN_2050; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_2051 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_33_out_out_out_7 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_3 = io_exe_rd_3_req_iscoef ? tmp_33_out_out_out_6 : tmp_33_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2056 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2057 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_2056; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2058 = 3'h3 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_2057; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2059 = 3'h4 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_2058; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_6 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2059 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2062 = 2'h1 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2063 = 2'h2 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_20_2 : _GEN_2062; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2064 = 2'h3 == _tmp_14_out_out_T_14[1:0] ? reg_type5_data_nxt_20_3 : _GEN_2063; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_7 = _tmp_14_out_out_T_14 < 3'h4 ? _GEN_2064 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_7 = io_exe_rd_3_req_isgroup ? tmp_34_out_out_out_7 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_3 = io_exe_rd_3_req_iscoef ? tmp_34_out_out_out_6 : tmp_34_out_out_7; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2069 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2070 = 3'h2 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2069; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2071 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2070; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2072 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2071; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2072 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_3 = io_exe_rd_3_req_iscoef ? tmp_35_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2076 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2077 = 3'h2 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2076; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2078 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2077; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2079 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2078; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2079 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_3 = io_exe_rd_3_req_iscoef ? tmp_36_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2083 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2084 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_2083; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2085 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2084; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2086 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2085; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2086 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_3 = io_exe_rd_3_req_iscoef ? tmp_37_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2090 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2091 = 3'h2 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2090; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2092 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2091; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2093 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2092; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2093 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_3 = io_exe_rd_3_req_iscoef ? tmp_38_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2097 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2098 = 3'h2 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2097; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2099 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2098; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2100 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2099; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2100 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_3 = io_exe_rd_3_req_iscoef ? tmp_39_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2104 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2105 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_2104; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2106 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2105; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2107 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2106; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2107 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_3 = io_exe_rd_3_req_iscoef ? tmp_40_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2111 = 3'h1 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2112 = 3'h2 == io_exe_rd_3_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_2111; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2113 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2112; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2114 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2113; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2114 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_3 = io_exe_rd_3_req_iscoef ? tmp_41_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2118 = 3'h1 == io_exe_rd_3_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2119 = 3'h2 == io_exe_rd_3_req_gidx ? reg_type6_coef_7_2 : _GEN_2118; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2120 = 3'h3 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2119; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2121 = 3'h4 == io_exe_rd_3_req_gidx ? 32'h0 : _GEN_2120; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_3 = io_exe_rd_3_req_gidx < 3'h5 ? _GEN_2121 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_3 = io_exe_rd_3_req_iscoef ? tmp_42_out_out_out_3 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_3 = io_exe_rd_3_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_3 = io_exe_rd_3_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_3 = io_exe_rd_3_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_3 = io_exe_rd_3_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_3 = io_exe_rd_3_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_3 = io_exe_rd_3_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_3 = io_exe_rd_3_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_3 = io_exe_rd_3_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_3_resp_T = 64'h1 << io_exe_rd_3_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_3_resp_T_52 = _io_exe_rd_3_resp_T[0] ? tmp_0_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_53 = _io_exe_rd_3_resp_T[1] ? tmp_1_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_54 = _io_exe_rd_3_resp_T[2] ? tmp_2_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_55 = _io_exe_rd_3_resp_T[3] ? tmp_3_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_56 = _io_exe_rd_3_resp_T[4] ? tmp_4_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_57 = _io_exe_rd_3_resp_T[5] ? tmp_5_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_58 = _io_exe_rd_3_resp_T[6] ? tmp_6_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_59 = _io_exe_rd_3_resp_T[7] ? tmp_7_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_60 = _io_exe_rd_3_resp_T[8] ? tmp_8_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_61 = _io_exe_rd_3_resp_T[9] ? tmp_9_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_62 = _io_exe_rd_3_resp_T[10] ? tmp_10_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_63 = _io_exe_rd_3_resp_T[11] ? tmp_11_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_64 = _io_exe_rd_3_resp_T[12] ? tmp_12_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_65 = _io_exe_rd_3_resp_T[13] ? tmp_13_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_66 = _io_exe_rd_3_resp_T[14] ? tmp_14_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_67 = _io_exe_rd_3_resp_T[15] ? tmp_15_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_68 = _io_exe_rd_3_resp_T[16] ? tmp_16_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_69 = _io_exe_rd_3_resp_T[17] ? tmp_17_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_70 = _io_exe_rd_3_resp_T[18] ? tmp_18_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_71 = _io_exe_rd_3_resp_T[19] ? tmp_19_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_72 = _io_exe_rd_3_resp_T[20] ? tmp_20_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_73 = _io_exe_rd_3_resp_T[21] ? tmp_21_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_74 = _io_exe_rd_3_resp_T[22] ? tmp_22_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_75 = _io_exe_rd_3_resp_T[23] ? tmp_23_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_76 = _io_exe_rd_3_resp_T[24] ? tmp_24_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_77 = _io_exe_rd_3_resp_T[25] ? tmp_25_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_78 = _io_exe_rd_3_resp_T[26] ? tmp_26_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_79 = _io_exe_rd_3_resp_T[27] ? tmp_27_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_80 = _io_exe_rd_3_resp_T[28] ? tmp_28_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_81 = _io_exe_rd_3_resp_T[29] ? tmp_29_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_82 = _io_exe_rd_3_resp_T[30] ? tmp_30_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_83 = _io_exe_rd_3_resp_T[31] ? tmp_31_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_84 = _io_exe_rd_3_resp_T[32] ? tmp_32_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_85 = _io_exe_rd_3_resp_T[33] ? tmp_33_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_86 = _io_exe_rd_3_resp_T[34] ? tmp_34_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_87 = _io_exe_rd_3_resp_T[35] ? tmp_35_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_88 = _io_exe_rd_3_resp_T[36] ? tmp_36_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_89 = _io_exe_rd_3_resp_T[37] ? tmp_37_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_90 = _io_exe_rd_3_resp_T[38] ? tmp_38_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_91 = _io_exe_rd_3_resp_T[39] ? tmp_39_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_92 = _io_exe_rd_3_resp_T[40] ? tmp_40_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_93 = _io_exe_rd_3_resp_T[41] ? tmp_41_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_94 = _io_exe_rd_3_resp_T[42] ? tmp_42_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_95 = _io_exe_rd_3_resp_T[43] ? tmp_43_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_96 = _io_exe_rd_3_resp_T[44] ? tmp_44_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_97 = _io_exe_rd_3_resp_T[45] ? tmp_45_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_98 = _io_exe_rd_3_resp_T[46] ? tmp_46_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_99 = _io_exe_rd_3_resp_T[47] ? tmp_47_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_100 = _io_exe_rd_3_resp_T[48] ? tmp_48_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_101 = _io_exe_rd_3_resp_T[49] ? tmp_49_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_102 = _io_exe_rd_3_resp_T[50] ? tmp_50_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_103 = _io_exe_rd_3_resp_T_52 | _io_exe_rd_3_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_104 = _io_exe_rd_3_resp_T_103 | _io_exe_rd_3_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_105 = _io_exe_rd_3_resp_T_104 | _io_exe_rd_3_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_106 = _io_exe_rd_3_resp_T_105 | _io_exe_rd_3_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_107 = _io_exe_rd_3_resp_T_106 | _io_exe_rd_3_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_108 = _io_exe_rd_3_resp_T_107 | _io_exe_rd_3_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_109 = _io_exe_rd_3_resp_T_108 | _io_exe_rd_3_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_110 = _io_exe_rd_3_resp_T_109 | _io_exe_rd_3_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_111 = _io_exe_rd_3_resp_T_110 | _io_exe_rd_3_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_112 = _io_exe_rd_3_resp_T_111 | _io_exe_rd_3_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_113 = _io_exe_rd_3_resp_T_112 | _io_exe_rd_3_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_114 = _io_exe_rd_3_resp_T_113 | _io_exe_rd_3_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_115 = _io_exe_rd_3_resp_T_114 | _io_exe_rd_3_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_116 = _io_exe_rd_3_resp_T_115 | _io_exe_rd_3_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_117 = _io_exe_rd_3_resp_T_116 | _io_exe_rd_3_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_118 = _io_exe_rd_3_resp_T_117 | _io_exe_rd_3_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_119 = _io_exe_rd_3_resp_T_118 | _io_exe_rd_3_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_120 = _io_exe_rd_3_resp_T_119 | _io_exe_rd_3_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_121 = _io_exe_rd_3_resp_T_120 | _io_exe_rd_3_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_122 = _io_exe_rd_3_resp_T_121 | _io_exe_rd_3_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_123 = _io_exe_rd_3_resp_T_122 | _io_exe_rd_3_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_124 = _io_exe_rd_3_resp_T_123 | _io_exe_rd_3_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_125 = _io_exe_rd_3_resp_T_124 | _io_exe_rd_3_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_126 = _io_exe_rd_3_resp_T_125 | _io_exe_rd_3_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_127 = _io_exe_rd_3_resp_T_126 | _io_exe_rd_3_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_128 = _io_exe_rd_3_resp_T_127 | _io_exe_rd_3_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_129 = _io_exe_rd_3_resp_T_128 | _io_exe_rd_3_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_130 = _io_exe_rd_3_resp_T_129 | _io_exe_rd_3_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_131 = _io_exe_rd_3_resp_T_130 | _io_exe_rd_3_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_132 = _io_exe_rd_3_resp_T_131 | _io_exe_rd_3_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_133 = _io_exe_rd_3_resp_T_132 | _io_exe_rd_3_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_134 = _io_exe_rd_3_resp_T_133 | _io_exe_rd_3_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_135 = _io_exe_rd_3_resp_T_134 | _io_exe_rd_3_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_136 = _io_exe_rd_3_resp_T_135 | _io_exe_rd_3_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_137 = _io_exe_rd_3_resp_T_136 | _io_exe_rd_3_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_138 = _io_exe_rd_3_resp_T_137 | _io_exe_rd_3_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_139 = _io_exe_rd_3_resp_T_138 | _io_exe_rd_3_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_140 = _io_exe_rd_3_resp_T_139 | _io_exe_rd_3_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_141 = _io_exe_rd_3_resp_T_140 | _io_exe_rd_3_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_142 = _io_exe_rd_3_resp_T_141 | _io_exe_rd_3_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_143 = _io_exe_rd_3_resp_T_142 | _io_exe_rd_3_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_144 = _io_exe_rd_3_resp_T_143 | _io_exe_rd_3_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_145 = _io_exe_rd_3_resp_T_144 | _io_exe_rd_3_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_146 = _io_exe_rd_3_resp_T_145 | _io_exe_rd_3_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_147 = _io_exe_rd_3_resp_T_146 | _io_exe_rd_3_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_148 = _io_exe_rd_3_resp_T_147 | _io_exe_rd_3_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_149 = _io_exe_rd_3_resp_T_148 | _io_exe_rd_3_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_150 = _io_exe_rd_3_resp_T_149 | _io_exe_rd_3_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_3_resp_T_151 = _io_exe_rd_3_resp_T_150 | _io_exe_rd_3_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_4 = io_exe_rd_4_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2141 = io_exe_rd_4_req_gidx[0] ? io_coef_in_mainch_drc_smooth_1 : io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h2 ? _GEN_2141 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_4 = io_exe_rd_4_req_iscoef ? tmp_8_out_out_out_4 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2145 = io_exe_rd_4_req_gidx[0] ? io_coef_in_subch_drc_smooth_1 : io_coef_in_subch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h2 ? _GEN_2145 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_4 = io_exe_rd_4_req_iscoef ? tmp_9_out_out_out_4 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2149 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2150 = 3'h2 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2149; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2151 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2150; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2152 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2151; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2152 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_4 = io_exe_rd_4_req_iscoef ? tmp_10_out_out_out_4 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_4 = io_exe_rd_4_req_iscoef ? tmp_10_out_out_out_4 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2163 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2164 = 3'h2 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2163; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2165 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2164; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2166 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2165; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2166 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_4 = io_exe_rd_4_req_iscoef ? tmp_12_out_out_out_4 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_4 = io_exe_rd_4_req_iscoef ? tmp_12_out_out_out_4 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2177 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2178 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_2177; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2179 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_2178; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2180 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_2179; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2180 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_18 = io_exe_rd_4_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_2183 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2184 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt__2 : _GEN_2183; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2185 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt__3 : _GEN_2184; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2185 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_14_out_out_out_9 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_4 = io_exe_rd_4_req_iscoef ? tmp_14_out_out_out_8 : tmp_14_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2190 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2191 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_2190; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2192 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_2191; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2193 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_2192; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2193 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2196 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2197 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_1_2 : _GEN_2196; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2198 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_1_3 : _GEN_2197; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2198 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_15_out_out_out_9 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_4 = io_exe_rd_4_req_iscoef ? tmp_15_out_out_out_8 : tmp_15_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2203 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2204 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_2203; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2205 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_2204; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2206 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_2205; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2206 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2209 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2210 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_2_2 : _GEN_2209; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2211 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_2_3 : _GEN_2210; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2211 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_16_out_out_out_9 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_4 = io_exe_rd_4_req_iscoef ? tmp_16_out_out_out_8 : tmp_16_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2216 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2217 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_2216; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2218 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_2217; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2219 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_2218; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2219 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2222 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2223 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_3_2 : _GEN_2222; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2224 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_3_3 : _GEN_2223; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2224 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_17_out_out_out_9 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_4 = io_exe_rd_4_req_iscoef ? tmp_17_out_out_out_8 : tmp_17_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2229 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2230 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_2229; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2231 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_2230; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2232 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_2231; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2232 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2235 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2236 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_4_2 : _GEN_2235; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2237 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_4_3 : _GEN_2236; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2237 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_18_out_out_out_9 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_4 = io_exe_rd_4_req_iscoef ? tmp_18_out_out_out_8 : tmp_18_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2242 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2243 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_2242; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2244 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_2243; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2245 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_2244; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2245 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2248 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2249 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_5_2 : _GEN_2248; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2250 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_5_3 : _GEN_2249; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2250 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_19_out_out_out_9 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_4 = io_exe_rd_4_req_iscoef ? tmp_19_out_out_out_8 : tmp_19_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2255 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2256 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_2255; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2257 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_2256; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2258 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_2257; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2258 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2261 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2262 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_6_2 : _GEN_2261; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2263 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_6_3 : _GEN_2262; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2263 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_20_out_out_out_9 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_4 = io_exe_rd_4_req_iscoef ? tmp_20_out_out_out_8 : tmp_20_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2268 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2269 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_2268; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2270 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_2269; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2271 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_2270; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2271 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2274 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2275 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_7_2 : _GEN_2274; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2276 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_7_3 : _GEN_2275; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2276 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_21_out_out_out_9 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_4 = io_exe_rd_4_req_iscoef ? tmp_21_out_out_out_8 : tmp_21_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2281 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2282 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_2281; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2283 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_2282; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2284 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_2283; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2284 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2287 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2288 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_8_2 : _GEN_2287; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2289 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_8_3 : _GEN_2288; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2289 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_22_out_out_out_9 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_4 = io_exe_rd_4_req_iscoef ? tmp_22_out_out_out_8 : tmp_22_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2294 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2295 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_2294; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2296 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_2295; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2297 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_2296; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2297 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2300 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2301 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_9_2 : _GEN_2300; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2302 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_9_3 : _GEN_2301; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2302 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_23_out_out_out_9 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_4 = io_exe_rd_4_req_iscoef ? tmp_23_out_out_out_8 : tmp_23_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2307 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2308 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_2307; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2309 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_2308; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2310 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_2309; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2310 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2313 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2314 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_10_2 : _GEN_2313; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2315 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_10_3 : _GEN_2314; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2315 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_24_out_out_out_9 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_4 = io_exe_rd_4_req_iscoef ? tmp_24_out_out_out_8 : tmp_24_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2320 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2321 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_2320; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2322 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_2321; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2323 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_2322; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2323 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2326 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2327 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_11_2 : _GEN_2326; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2328 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_11_3 : _GEN_2327; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2328 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_25_out_out_out_9 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_4 = io_exe_rd_4_req_iscoef ? tmp_25_out_out_out_8 : tmp_25_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2333 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2334 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_2333; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2335 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_2334; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2336 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_2335; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2336 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2339 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2340 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_12_2 : _GEN_2339; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2341 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_12_3 : _GEN_2340; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2341 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_26_out_out_out_9 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_4 = io_exe_rd_4_req_iscoef ? tmp_26_out_out_out_8 : tmp_26_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2346 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2347 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_2346; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2348 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_2347; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2349 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_2348; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2349 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2352 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2353 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_13_2 : _GEN_2352; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2354 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_13_3 : _GEN_2353; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2354 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_27_out_out_out_9 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_4 = io_exe_rd_4_req_iscoef ? tmp_27_out_out_out_8 : tmp_27_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2359 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2360 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_2359; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2361 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_2360; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2362 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_2361; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2362 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2365 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2366 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_14_2 : _GEN_2365; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2367 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_14_3 : _GEN_2366; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2367 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_28_out_out_out_9 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_4 = io_exe_rd_4_req_iscoef ? tmp_28_out_out_out_8 : tmp_28_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2372 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2373 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_2372; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2374 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_2373; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2375 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_2374; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2375 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2378 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2379 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_15_2 : _GEN_2378; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2380 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_15_3 : _GEN_2379; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2380 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_29_out_out_out_9 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_4 = io_exe_rd_4_req_iscoef ? tmp_29_out_out_out_8 : tmp_29_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2385 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2386 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_2385; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2387 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_2386; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2388 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_2387; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2388 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2391 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2392 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_16_2 : _GEN_2391; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2393 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_16_3 : _GEN_2392; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2393 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_30_out_out_out_9 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_4 = io_exe_rd_4_req_iscoef ? tmp_30_out_out_out_8 : tmp_30_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2398 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2399 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_2398; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2400 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_2399; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2401 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_2400; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2401 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2404 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2405 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_17_2 : _GEN_2404; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2406 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_17_3 : _GEN_2405; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2406 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_31_out_out_out_9 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_4 = io_exe_rd_4_req_iscoef ? tmp_31_out_out_out_8 : tmp_31_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2411 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2412 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_2411; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2413 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_2412; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2414 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_2413; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2414 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2417 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2418 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_18_2 : _GEN_2417; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2419 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_18_3 : _GEN_2418; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2419 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_32_out_out_out_9 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_4 = io_exe_rd_4_req_iscoef ? tmp_32_out_out_out_8 : tmp_32_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2424 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2425 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_2424; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2426 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_2425; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2427 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_2426; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2427 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2430 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2431 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_19_2 : _GEN_2430; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2432 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_19_3 : _GEN_2431; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2432 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_33_out_out_out_9 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_4 = io_exe_rd_4_req_iscoef ? tmp_33_out_out_out_8 : tmp_33_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2437 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2438 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_2437; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2439 = 3'h3 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_2438; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2440 = 3'h4 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_2439; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_8 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2440 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2443 = 2'h1 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2444 = 2'h2 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_20_2 : _GEN_2443; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2445 = 2'h3 == _tmp_14_out_out_T_18[1:0] ? reg_type5_data_nxt_20_3 : _GEN_2444; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_9 = _tmp_14_out_out_T_18 < 3'h4 ? _GEN_2445 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_9 = io_exe_rd_4_req_isgroup ? tmp_34_out_out_out_9 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_4 = io_exe_rd_4_req_iscoef ? tmp_34_out_out_out_8 : tmp_34_out_out_9; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2450 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2451 = 3'h2 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2450; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2452 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2451; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2453 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2452; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2453 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_4 = io_exe_rd_4_req_iscoef ? tmp_35_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2457 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2458 = 3'h2 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2457; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2459 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2458; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2460 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2459; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2460 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_4 = io_exe_rd_4_req_iscoef ? tmp_36_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2464 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2465 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_2464; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2466 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2465; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2467 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2466; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2467 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_4 = io_exe_rd_4_req_iscoef ? tmp_37_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2471 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2472 = 3'h2 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2471; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2473 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2472; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2474 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2473; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2474 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_4 = io_exe_rd_4_req_iscoef ? tmp_38_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2478 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2479 = 3'h2 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2478; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2480 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2479; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2481 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2480; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2481 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_4 = io_exe_rd_4_req_iscoef ? tmp_39_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2485 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2486 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_2485; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2487 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2486; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2488 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2487; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2488 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_4 = io_exe_rd_4_req_iscoef ? tmp_40_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2492 = 3'h1 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2493 = 3'h2 == io_exe_rd_4_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_2492; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2494 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2493; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2495 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2494; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2495 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_4 = io_exe_rd_4_req_iscoef ? tmp_41_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2499 = 3'h1 == io_exe_rd_4_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2500 = 3'h2 == io_exe_rd_4_req_gidx ? reg_type6_coef_7_2 : _GEN_2499; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2501 = 3'h3 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2500; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2502 = 3'h4 == io_exe_rd_4_req_gidx ? 32'h0 : _GEN_2501; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_4 = io_exe_rd_4_req_gidx < 3'h5 ? _GEN_2502 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_4 = io_exe_rd_4_req_iscoef ? tmp_42_out_out_out_4 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_4 = io_exe_rd_4_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_4 = io_exe_rd_4_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_4 = io_exe_rd_4_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_4 = io_exe_rd_4_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_4 = io_exe_rd_4_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_4 = io_exe_rd_4_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_4 = io_exe_rd_4_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_4 = io_exe_rd_4_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_4_resp_T = 64'h1 << io_exe_rd_4_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_4_resp_T_52 = _io_exe_rd_4_resp_T[0] ? tmp_0_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_53 = _io_exe_rd_4_resp_T[1] ? tmp_1_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_54 = _io_exe_rd_4_resp_T[2] ? tmp_2_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_55 = _io_exe_rd_4_resp_T[3] ? tmp_3_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_56 = _io_exe_rd_4_resp_T[4] ? tmp_4_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_57 = _io_exe_rd_4_resp_T[5] ? tmp_5_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_58 = _io_exe_rd_4_resp_T[6] ? tmp_6_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_59 = _io_exe_rd_4_resp_T[7] ? tmp_7_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_60 = _io_exe_rd_4_resp_T[8] ? tmp_8_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_61 = _io_exe_rd_4_resp_T[9] ? tmp_9_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_62 = _io_exe_rd_4_resp_T[10] ? tmp_10_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_63 = _io_exe_rd_4_resp_T[11] ? tmp_11_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_64 = _io_exe_rd_4_resp_T[12] ? tmp_12_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_65 = _io_exe_rd_4_resp_T[13] ? tmp_13_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_66 = _io_exe_rd_4_resp_T[14] ? tmp_14_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_67 = _io_exe_rd_4_resp_T[15] ? tmp_15_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_68 = _io_exe_rd_4_resp_T[16] ? tmp_16_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_69 = _io_exe_rd_4_resp_T[17] ? tmp_17_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_70 = _io_exe_rd_4_resp_T[18] ? tmp_18_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_71 = _io_exe_rd_4_resp_T[19] ? tmp_19_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_72 = _io_exe_rd_4_resp_T[20] ? tmp_20_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_73 = _io_exe_rd_4_resp_T[21] ? tmp_21_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_74 = _io_exe_rd_4_resp_T[22] ? tmp_22_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_75 = _io_exe_rd_4_resp_T[23] ? tmp_23_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_76 = _io_exe_rd_4_resp_T[24] ? tmp_24_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_77 = _io_exe_rd_4_resp_T[25] ? tmp_25_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_78 = _io_exe_rd_4_resp_T[26] ? tmp_26_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_79 = _io_exe_rd_4_resp_T[27] ? tmp_27_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_80 = _io_exe_rd_4_resp_T[28] ? tmp_28_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_81 = _io_exe_rd_4_resp_T[29] ? tmp_29_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_82 = _io_exe_rd_4_resp_T[30] ? tmp_30_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_83 = _io_exe_rd_4_resp_T[31] ? tmp_31_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_84 = _io_exe_rd_4_resp_T[32] ? tmp_32_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_85 = _io_exe_rd_4_resp_T[33] ? tmp_33_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_86 = _io_exe_rd_4_resp_T[34] ? tmp_34_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_87 = _io_exe_rd_4_resp_T[35] ? tmp_35_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_88 = _io_exe_rd_4_resp_T[36] ? tmp_36_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_89 = _io_exe_rd_4_resp_T[37] ? tmp_37_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_90 = _io_exe_rd_4_resp_T[38] ? tmp_38_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_91 = _io_exe_rd_4_resp_T[39] ? tmp_39_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_92 = _io_exe_rd_4_resp_T[40] ? tmp_40_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_93 = _io_exe_rd_4_resp_T[41] ? tmp_41_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_94 = _io_exe_rd_4_resp_T[42] ? tmp_42_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_95 = _io_exe_rd_4_resp_T[43] ? tmp_43_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_96 = _io_exe_rd_4_resp_T[44] ? tmp_44_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_97 = _io_exe_rd_4_resp_T[45] ? tmp_45_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_98 = _io_exe_rd_4_resp_T[46] ? tmp_46_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_99 = _io_exe_rd_4_resp_T[47] ? tmp_47_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_100 = _io_exe_rd_4_resp_T[48] ? tmp_48_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_101 = _io_exe_rd_4_resp_T[49] ? tmp_49_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_102 = _io_exe_rd_4_resp_T[50] ? tmp_50_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_103 = _io_exe_rd_4_resp_T_52 | _io_exe_rd_4_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_104 = _io_exe_rd_4_resp_T_103 | _io_exe_rd_4_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_105 = _io_exe_rd_4_resp_T_104 | _io_exe_rd_4_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_106 = _io_exe_rd_4_resp_T_105 | _io_exe_rd_4_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_107 = _io_exe_rd_4_resp_T_106 | _io_exe_rd_4_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_108 = _io_exe_rd_4_resp_T_107 | _io_exe_rd_4_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_109 = _io_exe_rd_4_resp_T_108 | _io_exe_rd_4_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_110 = _io_exe_rd_4_resp_T_109 | _io_exe_rd_4_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_111 = _io_exe_rd_4_resp_T_110 | _io_exe_rd_4_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_112 = _io_exe_rd_4_resp_T_111 | _io_exe_rd_4_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_113 = _io_exe_rd_4_resp_T_112 | _io_exe_rd_4_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_114 = _io_exe_rd_4_resp_T_113 | _io_exe_rd_4_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_115 = _io_exe_rd_4_resp_T_114 | _io_exe_rd_4_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_116 = _io_exe_rd_4_resp_T_115 | _io_exe_rd_4_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_117 = _io_exe_rd_4_resp_T_116 | _io_exe_rd_4_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_118 = _io_exe_rd_4_resp_T_117 | _io_exe_rd_4_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_119 = _io_exe_rd_4_resp_T_118 | _io_exe_rd_4_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_120 = _io_exe_rd_4_resp_T_119 | _io_exe_rd_4_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_121 = _io_exe_rd_4_resp_T_120 | _io_exe_rd_4_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_122 = _io_exe_rd_4_resp_T_121 | _io_exe_rd_4_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_123 = _io_exe_rd_4_resp_T_122 | _io_exe_rd_4_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_124 = _io_exe_rd_4_resp_T_123 | _io_exe_rd_4_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_125 = _io_exe_rd_4_resp_T_124 | _io_exe_rd_4_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_126 = _io_exe_rd_4_resp_T_125 | _io_exe_rd_4_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_127 = _io_exe_rd_4_resp_T_126 | _io_exe_rd_4_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_128 = _io_exe_rd_4_resp_T_127 | _io_exe_rd_4_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_129 = _io_exe_rd_4_resp_T_128 | _io_exe_rd_4_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_130 = _io_exe_rd_4_resp_T_129 | _io_exe_rd_4_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_131 = _io_exe_rd_4_resp_T_130 | _io_exe_rd_4_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_132 = _io_exe_rd_4_resp_T_131 | _io_exe_rd_4_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_133 = _io_exe_rd_4_resp_T_132 | _io_exe_rd_4_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_134 = _io_exe_rd_4_resp_T_133 | _io_exe_rd_4_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_135 = _io_exe_rd_4_resp_T_134 | _io_exe_rd_4_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_136 = _io_exe_rd_4_resp_T_135 | _io_exe_rd_4_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_137 = _io_exe_rd_4_resp_T_136 | _io_exe_rd_4_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_138 = _io_exe_rd_4_resp_T_137 | _io_exe_rd_4_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_139 = _io_exe_rd_4_resp_T_138 | _io_exe_rd_4_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_140 = _io_exe_rd_4_resp_T_139 | _io_exe_rd_4_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_141 = _io_exe_rd_4_resp_T_140 | _io_exe_rd_4_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_142 = _io_exe_rd_4_resp_T_141 | _io_exe_rd_4_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_143 = _io_exe_rd_4_resp_T_142 | _io_exe_rd_4_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_144 = _io_exe_rd_4_resp_T_143 | _io_exe_rd_4_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_145 = _io_exe_rd_4_resp_T_144 | _io_exe_rd_4_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_146 = _io_exe_rd_4_resp_T_145 | _io_exe_rd_4_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_147 = _io_exe_rd_4_resp_T_146 | _io_exe_rd_4_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_148 = _io_exe_rd_4_resp_T_147 | _io_exe_rd_4_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_149 = _io_exe_rd_4_resp_T_148 | _io_exe_rd_4_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_150 = _io_exe_rd_4_resp_T_149 | _io_exe_rd_4_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_4_resp_T_151 = _io_exe_rd_4_resp_T_150 | _io_exe_rd_4_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_5 = io_exe_rd_5_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_8_out_coef_out_5_0 = io_exe_rd_5_req_sel ? io_coef_in_mainch_drc_smooth_2 :
    io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_8_out_coef_out_5_1 = io_exe_rd_5_req_sel ? io_coef_in_mainch_drc_smooth_3 :
    io_coef_in_mainch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_2522 = io_exe_rd_5_req_gidx[0] ? tmp_8_out_coef_out_5_1 : tmp_8_out_coef_out_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h2 ? _GEN_2522 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_5 = io_exe_rd_5_req_iscoef ? tmp_8_out_out_out_5 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_9_out_coef_out_5_0 = io_exe_rd_5_req_sel ? io_coef_in_subch_drc_smooth_2 :
    io_coef_in_subch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_9_out_coef_out_5_1 = io_exe_rd_5_req_sel ? io_coef_in_subch_drc_smooth_3 :
    io_coef_in_subch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_2526 = io_exe_rd_5_req_gidx[0] ? tmp_9_out_coef_out_5_1 : tmp_9_out_coef_out_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h2 ? _GEN_2526 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_5 = io_exe_rd_5_req_iscoef ? tmp_9_out_out_out_5 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2530 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2531 = 3'h2 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2530; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2532 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2531; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2533 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2532; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2533 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_5 = io_exe_rd_5_req_iscoef ? tmp_10_out_out_out_5 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_5 = io_exe_rd_5_req_iscoef ? tmp_10_out_out_out_5 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2544 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2545 = 3'h2 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2544; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2546 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2545; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2547 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2546; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2547 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_5 = io_exe_rd_5_req_iscoef ? tmp_12_out_out_out_5 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_5 = io_exe_rd_5_req_iscoef ? tmp_12_out_out_out_5 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2558 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2559 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_2558; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2560 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_2559; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2561 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_2560; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2561 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_22 = io_exe_rd_5_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_2564 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2565 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt__2 : _GEN_2564; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2566 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt__3 : _GEN_2565; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2566 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_14_out_out_out_11 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_5 = io_exe_rd_5_req_iscoef ? tmp_14_out_out_out_10 : tmp_14_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2571 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2572 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_2571; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2573 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_2572; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2574 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_2573; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2574 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2577 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2578 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_1_2 : _GEN_2577; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2579 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_1_3 : _GEN_2578; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2579 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_15_out_out_out_11 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_5 = io_exe_rd_5_req_iscoef ? tmp_15_out_out_out_10 : tmp_15_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2584 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2585 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_2584; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2586 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_2585; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2587 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_2586; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2587 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2590 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2591 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_2_2 : _GEN_2590; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2592 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_2_3 : _GEN_2591; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2592 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_16_out_out_out_11 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_5 = io_exe_rd_5_req_iscoef ? tmp_16_out_out_out_10 : tmp_16_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2597 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2598 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_2597; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2599 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_2598; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2600 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_2599; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2600 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2603 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2604 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_3_2 : _GEN_2603; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2605 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_3_3 : _GEN_2604; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2605 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_17_out_out_out_11 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_5 = io_exe_rd_5_req_iscoef ? tmp_17_out_out_out_10 : tmp_17_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2610 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2611 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_2610; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2612 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_2611; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2613 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_2612; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2613 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2616 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2617 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_4_2 : _GEN_2616; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2618 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_4_3 : _GEN_2617; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2618 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_18_out_out_out_11 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_5 = io_exe_rd_5_req_iscoef ? tmp_18_out_out_out_10 : tmp_18_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2623 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2624 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_2623; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2625 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_2624; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2626 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_2625; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2626 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2629 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2630 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_5_2 : _GEN_2629; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2631 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_5_3 : _GEN_2630; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2631 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_19_out_out_out_11 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_5 = io_exe_rd_5_req_iscoef ? tmp_19_out_out_out_10 : tmp_19_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2636 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2637 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_2636; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2638 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_2637; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2639 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_2638; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2639 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2642 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2643 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_6_2 : _GEN_2642; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2644 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_6_3 : _GEN_2643; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2644 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_20_out_out_out_11 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_5 = io_exe_rd_5_req_iscoef ? tmp_20_out_out_out_10 : tmp_20_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2649 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2650 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_2649; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2651 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_2650; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2652 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_2651; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2652 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2655 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2656 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_7_2 : _GEN_2655; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2657 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_7_3 : _GEN_2656; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2657 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_21_out_out_out_11 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_5 = io_exe_rd_5_req_iscoef ? tmp_21_out_out_out_10 : tmp_21_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2662 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2663 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_2662; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2664 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_2663; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2665 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_2664; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2665 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2668 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2669 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_8_2 : _GEN_2668; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2670 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_8_3 : _GEN_2669; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2670 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_22_out_out_out_11 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_5 = io_exe_rd_5_req_iscoef ? tmp_22_out_out_out_10 : tmp_22_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2675 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2676 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_2675; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2677 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_2676; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2678 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_2677; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2678 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2681 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2682 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_9_2 : _GEN_2681; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2683 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_9_3 : _GEN_2682; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2683 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_23_out_out_out_11 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_5 = io_exe_rd_5_req_iscoef ? tmp_23_out_out_out_10 : tmp_23_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2688 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2689 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_2688; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2690 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_2689; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2691 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_2690; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2691 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2694 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2695 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_10_2 : _GEN_2694; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2696 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_10_3 : _GEN_2695; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2696 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_24_out_out_out_11 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_5 = io_exe_rd_5_req_iscoef ? tmp_24_out_out_out_10 : tmp_24_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2701 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2702 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_2701; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2703 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_2702; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2704 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_2703; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2704 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2707 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2708 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_11_2 : _GEN_2707; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2709 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_11_3 : _GEN_2708; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2709 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_25_out_out_out_11 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_5 = io_exe_rd_5_req_iscoef ? tmp_25_out_out_out_10 : tmp_25_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2714 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2715 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_2714; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2716 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_2715; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2717 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_2716; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2717 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2720 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2721 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_12_2 : _GEN_2720; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2722 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_12_3 : _GEN_2721; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2722 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_26_out_out_out_11 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_5 = io_exe_rd_5_req_iscoef ? tmp_26_out_out_out_10 : tmp_26_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2727 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2728 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_2727; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2729 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_2728; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2730 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_2729; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2730 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2733 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2734 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_13_2 : _GEN_2733; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2735 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_13_3 : _GEN_2734; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2735 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_27_out_out_out_11 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_5 = io_exe_rd_5_req_iscoef ? tmp_27_out_out_out_10 : tmp_27_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2740 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2741 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_2740; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2742 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_2741; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2743 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_2742; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2743 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2746 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2747 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_14_2 : _GEN_2746; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2748 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_14_3 : _GEN_2747; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2748 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_28_out_out_out_11 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_5 = io_exe_rd_5_req_iscoef ? tmp_28_out_out_out_10 : tmp_28_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2753 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2754 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_2753; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2755 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_2754; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2756 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_2755; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2756 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2759 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2760 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_15_2 : _GEN_2759; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2761 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_15_3 : _GEN_2760; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2761 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_29_out_out_out_11 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_5 = io_exe_rd_5_req_iscoef ? tmp_29_out_out_out_10 : tmp_29_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2766 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2767 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_2766; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2768 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_2767; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2769 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_2768; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2769 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2772 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2773 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_16_2 : _GEN_2772; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2774 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_16_3 : _GEN_2773; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2774 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_30_out_out_out_11 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_5 = io_exe_rd_5_req_iscoef ? tmp_30_out_out_out_10 : tmp_30_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2779 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2780 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_2779; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2781 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_2780; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2782 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_2781; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2782 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2785 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2786 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_17_2 : _GEN_2785; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2787 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_17_3 : _GEN_2786; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2787 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_31_out_out_out_11 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_5 = io_exe_rd_5_req_iscoef ? tmp_31_out_out_out_10 : tmp_31_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2792 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2793 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_2792; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2794 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_2793; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2795 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_2794; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2795 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2798 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2799 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_18_2 : _GEN_2798; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2800 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_18_3 : _GEN_2799; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2800 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_32_out_out_out_11 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_5 = io_exe_rd_5_req_iscoef ? tmp_32_out_out_out_10 : tmp_32_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2805 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2806 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_2805; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2807 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_2806; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2808 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_2807; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2808 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2811 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2812 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_19_2 : _GEN_2811; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2813 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_19_3 : _GEN_2812; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2813 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_33_out_out_out_11 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_5 = io_exe_rd_5_req_iscoef ? tmp_33_out_out_out_10 : tmp_33_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2818 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2819 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_2818; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2820 = 3'h3 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_2819; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2821 = 3'h4 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_2820; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_10 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2821 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2824 = 2'h1 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2825 = 2'h2 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_20_2 : _GEN_2824; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2826 = 2'h3 == _tmp_14_out_out_T_22[1:0] ? reg_type5_data_nxt_20_3 : _GEN_2825; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_11 = _tmp_14_out_out_T_22 < 3'h4 ? _GEN_2826 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_11 = io_exe_rd_5_req_isgroup ? tmp_34_out_out_out_11 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_5 = io_exe_rd_5_req_iscoef ? tmp_34_out_out_out_10 : tmp_34_out_out_11; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2831 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2832 = 3'h2 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2831; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2833 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2832; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2834 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2833; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2834 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_5 = io_exe_rd_5_req_iscoef ? tmp_35_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2838 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2839 = 3'h2 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2838; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2840 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2839; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2841 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2840; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2841 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_5 = io_exe_rd_5_req_iscoef ? tmp_36_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2845 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2846 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_2845; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2847 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2846; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2848 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2847; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2848 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_5 = io_exe_rd_5_req_iscoef ? tmp_37_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2852 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2853 = 3'h2 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2852; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2854 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2853; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2855 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2854; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2855 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_5 = io_exe_rd_5_req_iscoef ? tmp_38_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2859 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2860 = 3'h2 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2859; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2861 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2860; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2862 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2861; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2862 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_5 = io_exe_rd_5_req_iscoef ? tmp_39_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2866 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2867 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_2866; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2868 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2867; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2869 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2868; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2869 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_5 = io_exe_rd_5_req_iscoef ? tmp_40_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2873 = 3'h1 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2874 = 3'h2 == io_exe_rd_5_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_2873; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2875 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2874; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2876 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2875; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2876 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_5 = io_exe_rd_5_req_iscoef ? tmp_41_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2880 = 3'h1 == io_exe_rd_5_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2881 = 3'h2 == io_exe_rd_5_req_gidx ? reg_type6_coef_7_2 : _GEN_2880; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2882 = 3'h3 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2881; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2883 = 3'h4 == io_exe_rd_5_req_gidx ? 32'h0 : _GEN_2882; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_5 = io_exe_rd_5_req_gidx < 3'h5 ? _GEN_2883 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_5 = io_exe_rd_5_req_iscoef ? tmp_42_out_out_out_5 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_5 = io_exe_rd_5_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_5 = io_exe_rd_5_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_5 = io_exe_rd_5_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_5 = io_exe_rd_5_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_5 = io_exe_rd_5_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_5 = io_exe_rd_5_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_5 = io_exe_rd_5_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_5 = io_exe_rd_5_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_5_resp_T = 64'h1 << io_exe_rd_5_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_5_resp_T_52 = _io_exe_rd_5_resp_T[0] ? tmp_0_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_53 = _io_exe_rd_5_resp_T[1] ? tmp_1_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_54 = _io_exe_rd_5_resp_T[2] ? tmp_2_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_55 = _io_exe_rd_5_resp_T[3] ? tmp_3_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_56 = _io_exe_rd_5_resp_T[4] ? tmp_4_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_57 = _io_exe_rd_5_resp_T[5] ? tmp_5_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_58 = _io_exe_rd_5_resp_T[6] ? tmp_6_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_59 = _io_exe_rd_5_resp_T[7] ? tmp_7_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_60 = _io_exe_rd_5_resp_T[8] ? tmp_8_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_61 = _io_exe_rd_5_resp_T[9] ? tmp_9_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_62 = _io_exe_rd_5_resp_T[10] ? tmp_10_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_63 = _io_exe_rd_5_resp_T[11] ? tmp_11_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_64 = _io_exe_rd_5_resp_T[12] ? tmp_12_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_65 = _io_exe_rd_5_resp_T[13] ? tmp_13_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_66 = _io_exe_rd_5_resp_T[14] ? tmp_14_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_67 = _io_exe_rd_5_resp_T[15] ? tmp_15_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_68 = _io_exe_rd_5_resp_T[16] ? tmp_16_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_69 = _io_exe_rd_5_resp_T[17] ? tmp_17_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_70 = _io_exe_rd_5_resp_T[18] ? tmp_18_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_71 = _io_exe_rd_5_resp_T[19] ? tmp_19_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_72 = _io_exe_rd_5_resp_T[20] ? tmp_20_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_73 = _io_exe_rd_5_resp_T[21] ? tmp_21_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_74 = _io_exe_rd_5_resp_T[22] ? tmp_22_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_75 = _io_exe_rd_5_resp_T[23] ? tmp_23_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_76 = _io_exe_rd_5_resp_T[24] ? tmp_24_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_77 = _io_exe_rd_5_resp_T[25] ? tmp_25_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_78 = _io_exe_rd_5_resp_T[26] ? tmp_26_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_79 = _io_exe_rd_5_resp_T[27] ? tmp_27_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_80 = _io_exe_rd_5_resp_T[28] ? tmp_28_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_81 = _io_exe_rd_5_resp_T[29] ? tmp_29_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_82 = _io_exe_rd_5_resp_T[30] ? tmp_30_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_83 = _io_exe_rd_5_resp_T[31] ? tmp_31_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_84 = _io_exe_rd_5_resp_T[32] ? tmp_32_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_85 = _io_exe_rd_5_resp_T[33] ? tmp_33_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_86 = _io_exe_rd_5_resp_T[34] ? tmp_34_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_87 = _io_exe_rd_5_resp_T[35] ? tmp_35_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_88 = _io_exe_rd_5_resp_T[36] ? tmp_36_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_89 = _io_exe_rd_5_resp_T[37] ? tmp_37_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_90 = _io_exe_rd_5_resp_T[38] ? tmp_38_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_91 = _io_exe_rd_5_resp_T[39] ? tmp_39_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_92 = _io_exe_rd_5_resp_T[40] ? tmp_40_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_93 = _io_exe_rd_5_resp_T[41] ? tmp_41_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_94 = _io_exe_rd_5_resp_T[42] ? tmp_42_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_95 = _io_exe_rd_5_resp_T[43] ? tmp_43_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_96 = _io_exe_rd_5_resp_T[44] ? tmp_44_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_97 = _io_exe_rd_5_resp_T[45] ? tmp_45_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_98 = _io_exe_rd_5_resp_T[46] ? tmp_46_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_99 = _io_exe_rd_5_resp_T[47] ? tmp_47_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_100 = _io_exe_rd_5_resp_T[48] ? tmp_48_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_101 = _io_exe_rd_5_resp_T[49] ? tmp_49_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_102 = _io_exe_rd_5_resp_T[50] ? tmp_50_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_103 = _io_exe_rd_5_resp_T_52 | _io_exe_rd_5_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_104 = _io_exe_rd_5_resp_T_103 | _io_exe_rd_5_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_105 = _io_exe_rd_5_resp_T_104 | _io_exe_rd_5_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_106 = _io_exe_rd_5_resp_T_105 | _io_exe_rd_5_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_107 = _io_exe_rd_5_resp_T_106 | _io_exe_rd_5_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_108 = _io_exe_rd_5_resp_T_107 | _io_exe_rd_5_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_109 = _io_exe_rd_5_resp_T_108 | _io_exe_rd_5_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_110 = _io_exe_rd_5_resp_T_109 | _io_exe_rd_5_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_111 = _io_exe_rd_5_resp_T_110 | _io_exe_rd_5_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_112 = _io_exe_rd_5_resp_T_111 | _io_exe_rd_5_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_113 = _io_exe_rd_5_resp_T_112 | _io_exe_rd_5_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_114 = _io_exe_rd_5_resp_T_113 | _io_exe_rd_5_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_115 = _io_exe_rd_5_resp_T_114 | _io_exe_rd_5_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_116 = _io_exe_rd_5_resp_T_115 | _io_exe_rd_5_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_117 = _io_exe_rd_5_resp_T_116 | _io_exe_rd_5_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_118 = _io_exe_rd_5_resp_T_117 | _io_exe_rd_5_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_119 = _io_exe_rd_5_resp_T_118 | _io_exe_rd_5_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_120 = _io_exe_rd_5_resp_T_119 | _io_exe_rd_5_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_121 = _io_exe_rd_5_resp_T_120 | _io_exe_rd_5_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_122 = _io_exe_rd_5_resp_T_121 | _io_exe_rd_5_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_123 = _io_exe_rd_5_resp_T_122 | _io_exe_rd_5_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_124 = _io_exe_rd_5_resp_T_123 | _io_exe_rd_5_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_125 = _io_exe_rd_5_resp_T_124 | _io_exe_rd_5_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_126 = _io_exe_rd_5_resp_T_125 | _io_exe_rd_5_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_127 = _io_exe_rd_5_resp_T_126 | _io_exe_rd_5_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_128 = _io_exe_rd_5_resp_T_127 | _io_exe_rd_5_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_129 = _io_exe_rd_5_resp_T_128 | _io_exe_rd_5_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_130 = _io_exe_rd_5_resp_T_129 | _io_exe_rd_5_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_131 = _io_exe_rd_5_resp_T_130 | _io_exe_rd_5_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_132 = _io_exe_rd_5_resp_T_131 | _io_exe_rd_5_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_133 = _io_exe_rd_5_resp_T_132 | _io_exe_rd_5_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_134 = _io_exe_rd_5_resp_T_133 | _io_exe_rd_5_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_135 = _io_exe_rd_5_resp_T_134 | _io_exe_rd_5_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_136 = _io_exe_rd_5_resp_T_135 | _io_exe_rd_5_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_137 = _io_exe_rd_5_resp_T_136 | _io_exe_rd_5_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_138 = _io_exe_rd_5_resp_T_137 | _io_exe_rd_5_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_139 = _io_exe_rd_5_resp_T_138 | _io_exe_rd_5_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_140 = _io_exe_rd_5_resp_T_139 | _io_exe_rd_5_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_141 = _io_exe_rd_5_resp_T_140 | _io_exe_rd_5_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_142 = _io_exe_rd_5_resp_T_141 | _io_exe_rd_5_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_143 = _io_exe_rd_5_resp_T_142 | _io_exe_rd_5_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_144 = _io_exe_rd_5_resp_T_143 | _io_exe_rd_5_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_145 = _io_exe_rd_5_resp_T_144 | _io_exe_rd_5_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_146 = _io_exe_rd_5_resp_T_145 | _io_exe_rd_5_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_147 = _io_exe_rd_5_resp_T_146 | _io_exe_rd_5_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_148 = _io_exe_rd_5_resp_T_147 | _io_exe_rd_5_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_149 = _io_exe_rd_5_resp_T_148 | _io_exe_rd_5_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_150 = _io_exe_rd_5_resp_T_149 | _io_exe_rd_5_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_5_resp_T_151 = _io_exe_rd_5_resp_T_150 | _io_exe_rd_5_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_6 = io_exe_rd_6_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2903 = io_exe_rd_6_req_gidx[0] ? io_coef_in_mainch_drc_smooth_1 : io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h2 ? _GEN_2903 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_6 = io_exe_rd_6_req_iscoef ? tmp_8_out_out_out_6 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2907 = io_exe_rd_6_req_gidx[0] ? io_coef_in_subch_drc_smooth_1 : io_coef_in_subch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h2 ? _GEN_2907 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_6 = io_exe_rd_6_req_iscoef ? tmp_9_out_out_out_6 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2911 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2912 = 3'h2 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_2911; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2913 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_2912; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2914 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_2913; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2914 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_6 = io_exe_rd_6_req_iscoef ? tmp_10_out_out_out_6 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_6 = io_exe_rd_6_req_iscoef ? tmp_10_out_out_out_6 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2925 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2926 = 3'h2 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_2925; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2927 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_2926; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2928 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_2927; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2928 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_6 = io_exe_rd_6_req_iscoef ? tmp_12_out_out_out_6 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_6 = io_exe_rd_6_req_iscoef ? tmp_12_out_out_out_6 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2939 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2940 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_2939; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2941 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_2940; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2942 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_2941; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2942 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_26 = io_exe_rd_6_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_2945 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2946 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt__2 : _GEN_2945; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2947 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt__3 : _GEN_2946; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_2947 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_14_out_out_out_13 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_6 = io_exe_rd_6_req_iscoef ? tmp_14_out_out_out_12 : tmp_14_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2952 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2953 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_2952; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2954 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_2953; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2955 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_2954; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2955 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2958 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2959 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_1_2 : _GEN_2958; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2960 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_1_3 : _GEN_2959; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_2960 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_15_out_out_out_13 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_6 = io_exe_rd_6_req_iscoef ? tmp_15_out_out_out_12 : tmp_15_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2965 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2966 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_2965; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2967 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_2966; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2968 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_2967; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2968 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2971 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2972 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_2_2 : _GEN_2971; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2973 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_2_3 : _GEN_2972; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_2973 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_16_out_out_out_13 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_6 = io_exe_rd_6_req_iscoef ? tmp_16_out_out_out_12 : tmp_16_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2978 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2979 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_2978; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2980 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_2979; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2981 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_2980; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2981 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2984 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2985 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_3_2 : _GEN_2984; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2986 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_3_3 : _GEN_2985; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_2986 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_17_out_out_out_13 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_6 = io_exe_rd_6_req_iscoef ? tmp_17_out_out_out_12 : tmp_17_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_2991 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2992 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_2991; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2993 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_2992; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2994 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_2993; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_2994 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_2997 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2998 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_4_2 : _GEN_2997; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_2999 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_4_3 : _GEN_2998; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_2999 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_18_out_out_out_13 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_6 = io_exe_rd_6_req_iscoef ? tmp_18_out_out_out_12 : tmp_18_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3004 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3005 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_3004; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3006 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_3005; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3007 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_3006; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3007 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3010 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3011 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_5_2 : _GEN_3010; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3012 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_5_3 : _GEN_3011; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3012 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_19_out_out_out_13 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_6 = io_exe_rd_6_req_iscoef ? tmp_19_out_out_out_12 : tmp_19_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3017 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3018 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_3017; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3019 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_3018; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3020 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_3019; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3020 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3023 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3024 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_6_2 : _GEN_3023; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3025 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_6_3 : _GEN_3024; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3025 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_20_out_out_out_13 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_6 = io_exe_rd_6_req_iscoef ? tmp_20_out_out_out_12 : tmp_20_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3030 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3031 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_3030; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3032 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_3031; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3033 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_3032; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3033 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3036 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3037 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_7_2 : _GEN_3036; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3038 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_7_3 : _GEN_3037; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3038 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_21_out_out_out_13 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_6 = io_exe_rd_6_req_iscoef ? tmp_21_out_out_out_12 : tmp_21_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3043 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3044 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_3043; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3045 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_3044; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3046 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_3045; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3046 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3049 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3050 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_8_2 : _GEN_3049; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3051 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_8_3 : _GEN_3050; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3051 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_22_out_out_out_13 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_6 = io_exe_rd_6_req_iscoef ? tmp_22_out_out_out_12 : tmp_22_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3056 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3057 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_3056; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3058 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_3057; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3059 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_3058; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3059 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3062 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3063 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_9_2 : _GEN_3062; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3064 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_9_3 : _GEN_3063; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3064 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_23_out_out_out_13 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_6 = io_exe_rd_6_req_iscoef ? tmp_23_out_out_out_12 : tmp_23_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3069 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3070 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_3069; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3071 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_3070; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3072 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_3071; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3072 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3075 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3076 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_10_2 : _GEN_3075; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3077 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_10_3 : _GEN_3076; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3077 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_24_out_out_out_13 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_6 = io_exe_rd_6_req_iscoef ? tmp_24_out_out_out_12 : tmp_24_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3082 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3083 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_3082; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3084 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_3083; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3085 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_3084; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3085 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3088 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3089 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_11_2 : _GEN_3088; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3090 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_11_3 : _GEN_3089; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3090 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_25_out_out_out_13 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_6 = io_exe_rd_6_req_iscoef ? tmp_25_out_out_out_12 : tmp_25_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3095 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3096 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_3095; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3097 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_3096; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3098 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_3097; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3098 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3101 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3102 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_12_2 : _GEN_3101; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3103 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_12_3 : _GEN_3102; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3103 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_26_out_out_out_13 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_6 = io_exe_rd_6_req_iscoef ? tmp_26_out_out_out_12 : tmp_26_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3108 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3109 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_3108; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3110 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_3109; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3111 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_3110; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3111 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3114 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3115 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_13_2 : _GEN_3114; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3116 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_13_3 : _GEN_3115; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3116 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_27_out_out_out_13 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_6 = io_exe_rd_6_req_iscoef ? tmp_27_out_out_out_12 : tmp_27_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3121 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3122 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_3121; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3123 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_3122; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3124 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_3123; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3124 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3127 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3128 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_14_2 : _GEN_3127; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3129 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_14_3 : _GEN_3128; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3129 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_28_out_out_out_13 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_6 = io_exe_rd_6_req_iscoef ? tmp_28_out_out_out_12 : tmp_28_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3134 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3135 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_3134; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3136 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_3135; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3137 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_3136; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3137 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3140 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3141 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_15_2 : _GEN_3140; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3142 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_15_3 : _GEN_3141; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3142 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_29_out_out_out_13 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_6 = io_exe_rd_6_req_iscoef ? tmp_29_out_out_out_12 : tmp_29_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3147 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3148 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_3147; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3149 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_3148; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3150 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_3149; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3150 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3153 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3154 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_16_2 : _GEN_3153; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3155 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_16_3 : _GEN_3154; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3155 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_30_out_out_out_13 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_6 = io_exe_rd_6_req_iscoef ? tmp_30_out_out_out_12 : tmp_30_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3160 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3161 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_3160; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3162 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_3161; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3163 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_3162; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3163 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3166 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3167 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_17_2 : _GEN_3166; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3168 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_17_3 : _GEN_3167; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3168 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_31_out_out_out_13 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_6 = io_exe_rd_6_req_iscoef ? tmp_31_out_out_out_12 : tmp_31_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3173 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3174 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_3173; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3175 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_3174; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3176 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_3175; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3176 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3179 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3180 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_18_2 : _GEN_3179; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3181 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_18_3 : _GEN_3180; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3181 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_32_out_out_out_13 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_6 = io_exe_rd_6_req_iscoef ? tmp_32_out_out_out_12 : tmp_32_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3186 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3187 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_3186; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3188 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_3187; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3189 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_3188; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3189 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3192 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3193 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_19_2 : _GEN_3192; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3194 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_19_3 : _GEN_3193; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3194 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_33_out_out_out_13 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_6 = io_exe_rd_6_req_iscoef ? tmp_33_out_out_out_12 : tmp_33_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3199 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3200 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_3199; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3201 = 3'h3 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_3200; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3202 = 3'h4 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_3201; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_12 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3202 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3205 = 2'h1 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3206 = 2'h2 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_20_2 : _GEN_3205; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3207 = 2'h3 == _tmp_14_out_out_T_26[1:0] ? reg_type5_data_nxt_20_3 : _GEN_3206; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_13 = _tmp_14_out_out_T_26 < 3'h4 ? _GEN_3207 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_13 = io_exe_rd_6_req_isgroup ? tmp_34_out_out_out_13 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_6 = io_exe_rd_6_req_iscoef ? tmp_34_out_out_out_12 : tmp_34_out_out_13; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3212 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3213 = 3'h2 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3212; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3214 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3213; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3215 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3214; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3215 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_6 = io_exe_rd_6_req_iscoef ? tmp_35_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3219 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3220 = 3'h2 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3219; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3221 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3220; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3222 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3221; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3222 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_6 = io_exe_rd_6_req_iscoef ? tmp_36_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3226 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3227 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_3226; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3228 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3227; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3229 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3228; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3229 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_6 = io_exe_rd_6_req_iscoef ? tmp_37_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3233 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3234 = 3'h2 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3233; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3235 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3234; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3236 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3235; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3236 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_6 = io_exe_rd_6_req_iscoef ? tmp_38_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3240 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3241 = 3'h2 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3240; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3242 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3241; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3243 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3242; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3243 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_6 = io_exe_rd_6_req_iscoef ? tmp_39_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3247 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3248 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_3247; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3249 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3248; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3250 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3249; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3250 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_6 = io_exe_rd_6_req_iscoef ? tmp_40_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3254 = 3'h1 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3255 = 3'h2 == io_exe_rd_6_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_3254; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3256 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3255; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3257 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3256; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3257 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_6 = io_exe_rd_6_req_iscoef ? tmp_41_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3261 = 3'h1 == io_exe_rd_6_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3262 = 3'h2 == io_exe_rd_6_req_gidx ? reg_type6_coef_7_2 : _GEN_3261; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3263 = 3'h3 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3262; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3264 = 3'h4 == io_exe_rd_6_req_gidx ? 32'h0 : _GEN_3263; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_6 = io_exe_rd_6_req_gidx < 3'h5 ? _GEN_3264 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_6 = io_exe_rd_6_req_iscoef ? tmp_42_out_out_out_6 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_6 = io_exe_rd_6_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_6 = io_exe_rd_6_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_6 = io_exe_rd_6_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_6 = io_exe_rd_6_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_6 = io_exe_rd_6_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_6 = io_exe_rd_6_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_6 = io_exe_rd_6_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_6 = io_exe_rd_6_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_6_resp_T = 64'h1 << io_exe_rd_6_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_6_resp_T_52 = _io_exe_rd_6_resp_T[0] ? tmp_0_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_53 = _io_exe_rd_6_resp_T[1] ? tmp_1_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_54 = _io_exe_rd_6_resp_T[2] ? tmp_2_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_55 = _io_exe_rd_6_resp_T[3] ? tmp_3_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_56 = _io_exe_rd_6_resp_T[4] ? tmp_4_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_57 = _io_exe_rd_6_resp_T[5] ? tmp_5_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_58 = _io_exe_rd_6_resp_T[6] ? tmp_6_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_59 = _io_exe_rd_6_resp_T[7] ? tmp_7_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_60 = _io_exe_rd_6_resp_T[8] ? tmp_8_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_61 = _io_exe_rd_6_resp_T[9] ? tmp_9_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_62 = _io_exe_rd_6_resp_T[10] ? tmp_10_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_63 = _io_exe_rd_6_resp_T[11] ? tmp_11_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_64 = _io_exe_rd_6_resp_T[12] ? tmp_12_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_65 = _io_exe_rd_6_resp_T[13] ? tmp_13_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_66 = _io_exe_rd_6_resp_T[14] ? tmp_14_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_67 = _io_exe_rd_6_resp_T[15] ? tmp_15_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_68 = _io_exe_rd_6_resp_T[16] ? tmp_16_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_69 = _io_exe_rd_6_resp_T[17] ? tmp_17_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_70 = _io_exe_rd_6_resp_T[18] ? tmp_18_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_71 = _io_exe_rd_6_resp_T[19] ? tmp_19_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_72 = _io_exe_rd_6_resp_T[20] ? tmp_20_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_73 = _io_exe_rd_6_resp_T[21] ? tmp_21_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_74 = _io_exe_rd_6_resp_T[22] ? tmp_22_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_75 = _io_exe_rd_6_resp_T[23] ? tmp_23_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_76 = _io_exe_rd_6_resp_T[24] ? tmp_24_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_77 = _io_exe_rd_6_resp_T[25] ? tmp_25_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_78 = _io_exe_rd_6_resp_T[26] ? tmp_26_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_79 = _io_exe_rd_6_resp_T[27] ? tmp_27_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_80 = _io_exe_rd_6_resp_T[28] ? tmp_28_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_81 = _io_exe_rd_6_resp_T[29] ? tmp_29_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_82 = _io_exe_rd_6_resp_T[30] ? tmp_30_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_83 = _io_exe_rd_6_resp_T[31] ? tmp_31_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_84 = _io_exe_rd_6_resp_T[32] ? tmp_32_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_85 = _io_exe_rd_6_resp_T[33] ? tmp_33_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_86 = _io_exe_rd_6_resp_T[34] ? tmp_34_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_87 = _io_exe_rd_6_resp_T[35] ? tmp_35_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_88 = _io_exe_rd_6_resp_T[36] ? tmp_36_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_89 = _io_exe_rd_6_resp_T[37] ? tmp_37_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_90 = _io_exe_rd_6_resp_T[38] ? tmp_38_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_91 = _io_exe_rd_6_resp_T[39] ? tmp_39_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_92 = _io_exe_rd_6_resp_T[40] ? tmp_40_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_93 = _io_exe_rd_6_resp_T[41] ? tmp_41_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_94 = _io_exe_rd_6_resp_T[42] ? tmp_42_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_95 = _io_exe_rd_6_resp_T[43] ? tmp_43_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_96 = _io_exe_rd_6_resp_T[44] ? tmp_44_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_97 = _io_exe_rd_6_resp_T[45] ? tmp_45_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_98 = _io_exe_rd_6_resp_T[46] ? tmp_46_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_99 = _io_exe_rd_6_resp_T[47] ? tmp_47_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_100 = _io_exe_rd_6_resp_T[48] ? tmp_48_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_101 = _io_exe_rd_6_resp_T[49] ? tmp_49_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_102 = _io_exe_rd_6_resp_T[50] ? tmp_50_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_103 = _io_exe_rd_6_resp_T_52 | _io_exe_rd_6_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_104 = _io_exe_rd_6_resp_T_103 | _io_exe_rd_6_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_105 = _io_exe_rd_6_resp_T_104 | _io_exe_rd_6_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_106 = _io_exe_rd_6_resp_T_105 | _io_exe_rd_6_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_107 = _io_exe_rd_6_resp_T_106 | _io_exe_rd_6_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_108 = _io_exe_rd_6_resp_T_107 | _io_exe_rd_6_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_109 = _io_exe_rd_6_resp_T_108 | _io_exe_rd_6_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_110 = _io_exe_rd_6_resp_T_109 | _io_exe_rd_6_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_111 = _io_exe_rd_6_resp_T_110 | _io_exe_rd_6_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_112 = _io_exe_rd_6_resp_T_111 | _io_exe_rd_6_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_113 = _io_exe_rd_6_resp_T_112 | _io_exe_rd_6_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_114 = _io_exe_rd_6_resp_T_113 | _io_exe_rd_6_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_115 = _io_exe_rd_6_resp_T_114 | _io_exe_rd_6_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_116 = _io_exe_rd_6_resp_T_115 | _io_exe_rd_6_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_117 = _io_exe_rd_6_resp_T_116 | _io_exe_rd_6_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_118 = _io_exe_rd_6_resp_T_117 | _io_exe_rd_6_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_119 = _io_exe_rd_6_resp_T_118 | _io_exe_rd_6_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_120 = _io_exe_rd_6_resp_T_119 | _io_exe_rd_6_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_121 = _io_exe_rd_6_resp_T_120 | _io_exe_rd_6_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_122 = _io_exe_rd_6_resp_T_121 | _io_exe_rd_6_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_123 = _io_exe_rd_6_resp_T_122 | _io_exe_rd_6_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_124 = _io_exe_rd_6_resp_T_123 | _io_exe_rd_6_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_125 = _io_exe_rd_6_resp_T_124 | _io_exe_rd_6_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_126 = _io_exe_rd_6_resp_T_125 | _io_exe_rd_6_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_127 = _io_exe_rd_6_resp_T_126 | _io_exe_rd_6_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_128 = _io_exe_rd_6_resp_T_127 | _io_exe_rd_6_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_129 = _io_exe_rd_6_resp_T_128 | _io_exe_rd_6_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_130 = _io_exe_rd_6_resp_T_129 | _io_exe_rd_6_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_131 = _io_exe_rd_6_resp_T_130 | _io_exe_rd_6_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_132 = _io_exe_rd_6_resp_T_131 | _io_exe_rd_6_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_133 = _io_exe_rd_6_resp_T_132 | _io_exe_rd_6_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_134 = _io_exe_rd_6_resp_T_133 | _io_exe_rd_6_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_135 = _io_exe_rd_6_resp_T_134 | _io_exe_rd_6_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_136 = _io_exe_rd_6_resp_T_135 | _io_exe_rd_6_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_137 = _io_exe_rd_6_resp_T_136 | _io_exe_rd_6_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_138 = _io_exe_rd_6_resp_T_137 | _io_exe_rd_6_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_139 = _io_exe_rd_6_resp_T_138 | _io_exe_rd_6_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_140 = _io_exe_rd_6_resp_T_139 | _io_exe_rd_6_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_141 = _io_exe_rd_6_resp_T_140 | _io_exe_rd_6_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_142 = _io_exe_rd_6_resp_T_141 | _io_exe_rd_6_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_143 = _io_exe_rd_6_resp_T_142 | _io_exe_rd_6_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_144 = _io_exe_rd_6_resp_T_143 | _io_exe_rd_6_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_145 = _io_exe_rd_6_resp_T_144 | _io_exe_rd_6_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_146 = _io_exe_rd_6_resp_T_145 | _io_exe_rd_6_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_147 = _io_exe_rd_6_resp_T_146 | _io_exe_rd_6_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_148 = _io_exe_rd_6_resp_T_147 | _io_exe_rd_6_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_149 = _io_exe_rd_6_resp_T_148 | _io_exe_rd_6_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_150 = _io_exe_rd_6_resp_T_149 | _io_exe_rd_6_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_6_resp_T_151 = _io_exe_rd_6_resp_T_150 | _io_exe_rd_6_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_7 = io_exe_rd_7_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_8_out_coef_out_7_0 = io_exe_rd_7_req_sel ? io_coef_in_mainch_drc_smooth_2 :
    io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_8_out_coef_out_7_1 = io_exe_rd_7_req_sel ? io_coef_in_mainch_drc_smooth_3 :
    io_coef_in_mainch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_3284 = io_exe_rd_7_req_gidx[0] ? tmp_8_out_coef_out_7_1 : tmp_8_out_coef_out_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h2 ? _GEN_3284 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_7 = io_exe_rd_7_req_iscoef ? tmp_8_out_out_out_7 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_9_out_coef_out_7_0 = io_exe_rd_7_req_sel ? io_coef_in_subch_drc_smooth_2 :
    io_coef_in_subch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_9_out_coef_out_7_1 = io_exe_rd_7_req_sel ? io_coef_in_subch_drc_smooth_3 :
    io_coef_in_subch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_3288 = io_exe_rd_7_req_gidx[0] ? tmp_9_out_coef_out_7_1 : tmp_9_out_coef_out_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h2 ? _GEN_3288 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_7 = io_exe_rd_7_req_iscoef ? tmp_9_out_out_out_7 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3292 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3293 = 3'h2 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3292; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3294 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3293; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3295 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3294; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3295 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_7 = io_exe_rd_7_req_iscoef ? tmp_10_out_out_out_7 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_7 = io_exe_rd_7_req_iscoef ? tmp_10_out_out_out_7 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3306 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3307 = 3'h2 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3306; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3308 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3307; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3309 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3308; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3309 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_7 = io_exe_rd_7_req_iscoef ? tmp_12_out_out_out_7 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_7 = io_exe_rd_7_req_iscoef ? tmp_12_out_out_out_7 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3320 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3321 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_3320; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3322 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_3321; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3323 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_3322; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3323 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_30 = io_exe_rd_7_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_3326 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3327 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt__2 : _GEN_3326; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3328 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt__3 : _GEN_3327; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3328 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_14_out_out_out_15 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_7 = io_exe_rd_7_req_iscoef ? tmp_14_out_out_out_14 : tmp_14_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3333 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3334 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_3333; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3335 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_3334; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3336 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_3335; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3336 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3339 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3340 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_1_2 : _GEN_3339; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3341 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_1_3 : _GEN_3340; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3341 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_15_out_out_out_15 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_7 = io_exe_rd_7_req_iscoef ? tmp_15_out_out_out_14 : tmp_15_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3346 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3347 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_3346; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3348 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_3347; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3349 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_3348; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3349 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3352 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3353 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_2_2 : _GEN_3352; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3354 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_2_3 : _GEN_3353; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3354 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_16_out_out_out_15 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_7 = io_exe_rd_7_req_iscoef ? tmp_16_out_out_out_14 : tmp_16_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3359 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3360 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_3359; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3361 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_3360; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3362 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_3361; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3362 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3365 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3366 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_3_2 : _GEN_3365; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3367 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_3_3 : _GEN_3366; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3367 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_17_out_out_out_15 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_7 = io_exe_rd_7_req_iscoef ? tmp_17_out_out_out_14 : tmp_17_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3372 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3373 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_3372; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3374 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_3373; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3375 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_3374; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3375 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3378 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3379 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_4_2 : _GEN_3378; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3380 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_4_3 : _GEN_3379; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3380 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_18_out_out_out_15 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_7 = io_exe_rd_7_req_iscoef ? tmp_18_out_out_out_14 : tmp_18_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3385 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3386 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_3385; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3387 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_3386; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3388 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_3387; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3388 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3391 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3392 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_5_2 : _GEN_3391; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3393 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_5_3 : _GEN_3392; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3393 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_19_out_out_out_15 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_7 = io_exe_rd_7_req_iscoef ? tmp_19_out_out_out_14 : tmp_19_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3398 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3399 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_3398; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3400 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_3399; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3401 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_3400; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3401 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3404 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3405 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_6_2 : _GEN_3404; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3406 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_6_3 : _GEN_3405; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3406 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_20_out_out_out_15 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_7 = io_exe_rd_7_req_iscoef ? tmp_20_out_out_out_14 : tmp_20_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3411 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3412 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_3411; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3413 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_3412; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3414 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_3413; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3414 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3417 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3418 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_7_2 : _GEN_3417; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3419 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_7_3 : _GEN_3418; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3419 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_21_out_out_out_15 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_7 = io_exe_rd_7_req_iscoef ? tmp_21_out_out_out_14 : tmp_21_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3424 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3425 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_3424; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3426 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_3425; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3427 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_3426; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3427 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3430 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3431 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_8_2 : _GEN_3430; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3432 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_8_3 : _GEN_3431; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3432 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_22_out_out_out_15 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_7 = io_exe_rd_7_req_iscoef ? tmp_22_out_out_out_14 : tmp_22_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3437 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3438 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_3437; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3439 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_3438; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3440 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_3439; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3440 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3443 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3444 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_9_2 : _GEN_3443; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3445 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_9_3 : _GEN_3444; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3445 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_23_out_out_out_15 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_7 = io_exe_rd_7_req_iscoef ? tmp_23_out_out_out_14 : tmp_23_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3450 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3451 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_3450; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3452 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_3451; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3453 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_3452; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3453 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3456 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3457 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_10_2 : _GEN_3456; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3458 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_10_3 : _GEN_3457; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3458 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_24_out_out_out_15 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_7 = io_exe_rd_7_req_iscoef ? tmp_24_out_out_out_14 : tmp_24_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3463 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3464 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_3463; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3465 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_3464; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3466 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_3465; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3466 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3469 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3470 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_11_2 : _GEN_3469; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3471 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_11_3 : _GEN_3470; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3471 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_25_out_out_out_15 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_7 = io_exe_rd_7_req_iscoef ? tmp_25_out_out_out_14 : tmp_25_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3476 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3477 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_3476; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3478 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_3477; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3479 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_3478; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3479 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3482 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3483 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_12_2 : _GEN_3482; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3484 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_12_3 : _GEN_3483; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3484 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_26_out_out_out_15 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_7 = io_exe_rd_7_req_iscoef ? tmp_26_out_out_out_14 : tmp_26_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3489 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3490 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_3489; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3491 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_3490; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3492 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_3491; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3492 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3495 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3496 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_13_2 : _GEN_3495; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3497 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_13_3 : _GEN_3496; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3497 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_27_out_out_out_15 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_7 = io_exe_rd_7_req_iscoef ? tmp_27_out_out_out_14 : tmp_27_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3502 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3503 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_3502; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3504 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_3503; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3505 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_3504; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3505 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3508 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3509 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_14_2 : _GEN_3508; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3510 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_14_3 : _GEN_3509; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3510 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_28_out_out_out_15 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_7 = io_exe_rd_7_req_iscoef ? tmp_28_out_out_out_14 : tmp_28_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3515 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3516 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_3515; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3517 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_3516; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3518 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_3517; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3518 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3521 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3522 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_15_2 : _GEN_3521; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3523 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_15_3 : _GEN_3522; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3523 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_29_out_out_out_15 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_7 = io_exe_rd_7_req_iscoef ? tmp_29_out_out_out_14 : tmp_29_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3528 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3529 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_3528; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3530 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_3529; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3531 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_3530; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3531 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3534 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3535 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_16_2 : _GEN_3534; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3536 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_16_3 : _GEN_3535; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3536 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_30_out_out_out_15 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_7 = io_exe_rd_7_req_iscoef ? tmp_30_out_out_out_14 : tmp_30_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3541 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3542 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_3541; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3543 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_3542; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3544 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_3543; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3544 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3547 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3548 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_17_2 : _GEN_3547; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3549 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_17_3 : _GEN_3548; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3549 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_31_out_out_out_15 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_7 = io_exe_rd_7_req_iscoef ? tmp_31_out_out_out_14 : tmp_31_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3554 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3555 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_3554; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3556 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_3555; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3557 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_3556; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3557 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3560 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3561 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_18_2 : _GEN_3560; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3562 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_18_3 : _GEN_3561; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3562 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_32_out_out_out_15 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_7 = io_exe_rd_7_req_iscoef ? tmp_32_out_out_out_14 : tmp_32_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3567 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3568 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_3567; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3569 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_3568; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3570 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_3569; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3570 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3573 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3574 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_19_2 : _GEN_3573; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3575 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_19_3 : _GEN_3574; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3575 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_33_out_out_out_15 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_7 = io_exe_rd_7_req_iscoef ? tmp_33_out_out_out_14 : tmp_33_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3580 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3581 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_3580; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3582 = 3'h3 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_3581; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3583 = 3'h4 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_3582; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_14 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3583 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3586 = 2'h1 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3587 = 2'h2 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_20_2 : _GEN_3586; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3588 = 2'h3 == _tmp_14_out_out_T_30[1:0] ? reg_type5_data_nxt_20_3 : _GEN_3587; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_15 = _tmp_14_out_out_T_30 < 3'h4 ? _GEN_3588 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_15 = io_exe_rd_7_req_isgroup ? tmp_34_out_out_out_15 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_7 = io_exe_rd_7_req_iscoef ? tmp_34_out_out_out_14 : tmp_34_out_out_15; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3593 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3594 = 3'h2 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3593; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3595 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3594; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3596 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3595; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3596 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_7 = io_exe_rd_7_req_iscoef ? tmp_35_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3600 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3601 = 3'h2 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3600; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3602 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3601; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3603 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3602; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3603 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_7 = io_exe_rd_7_req_iscoef ? tmp_36_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3607 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3608 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_3607; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3609 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3608; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3610 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3609; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3610 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_7 = io_exe_rd_7_req_iscoef ? tmp_37_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3614 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3615 = 3'h2 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3614; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3616 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3615; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3617 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3616; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3617 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_7 = io_exe_rd_7_req_iscoef ? tmp_38_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3621 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3622 = 3'h2 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3621; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3623 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3622; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3624 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3623; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3624 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_7 = io_exe_rd_7_req_iscoef ? tmp_39_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3628 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3629 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_3628; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3630 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3629; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3631 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3630; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3631 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_7 = io_exe_rd_7_req_iscoef ? tmp_40_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3635 = 3'h1 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3636 = 3'h2 == io_exe_rd_7_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_3635; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3637 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3636; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3638 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3637; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3638 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_7 = io_exe_rd_7_req_iscoef ? tmp_41_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3642 = 3'h1 == io_exe_rd_7_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3643 = 3'h2 == io_exe_rd_7_req_gidx ? reg_type6_coef_7_2 : _GEN_3642; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3644 = 3'h3 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3643; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3645 = 3'h4 == io_exe_rd_7_req_gidx ? 32'h0 : _GEN_3644; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_7 = io_exe_rd_7_req_gidx < 3'h5 ? _GEN_3645 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_7 = io_exe_rd_7_req_iscoef ? tmp_42_out_out_out_7 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_7 = io_exe_rd_7_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_7 = io_exe_rd_7_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_7 = io_exe_rd_7_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_7 = io_exe_rd_7_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_7 = io_exe_rd_7_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_7 = io_exe_rd_7_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_7 = io_exe_rd_7_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_7 = io_exe_rd_7_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_7_resp_T = 64'h1 << io_exe_rd_7_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_7_resp_T_52 = _io_exe_rd_7_resp_T[0] ? tmp_0_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_53 = _io_exe_rd_7_resp_T[1] ? tmp_1_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_54 = _io_exe_rd_7_resp_T[2] ? tmp_2_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_55 = _io_exe_rd_7_resp_T[3] ? tmp_3_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_56 = _io_exe_rd_7_resp_T[4] ? tmp_4_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_57 = _io_exe_rd_7_resp_T[5] ? tmp_5_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_58 = _io_exe_rd_7_resp_T[6] ? tmp_6_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_59 = _io_exe_rd_7_resp_T[7] ? tmp_7_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_60 = _io_exe_rd_7_resp_T[8] ? tmp_8_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_61 = _io_exe_rd_7_resp_T[9] ? tmp_9_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_62 = _io_exe_rd_7_resp_T[10] ? tmp_10_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_63 = _io_exe_rd_7_resp_T[11] ? tmp_11_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_64 = _io_exe_rd_7_resp_T[12] ? tmp_12_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_65 = _io_exe_rd_7_resp_T[13] ? tmp_13_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_66 = _io_exe_rd_7_resp_T[14] ? tmp_14_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_67 = _io_exe_rd_7_resp_T[15] ? tmp_15_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_68 = _io_exe_rd_7_resp_T[16] ? tmp_16_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_69 = _io_exe_rd_7_resp_T[17] ? tmp_17_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_70 = _io_exe_rd_7_resp_T[18] ? tmp_18_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_71 = _io_exe_rd_7_resp_T[19] ? tmp_19_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_72 = _io_exe_rd_7_resp_T[20] ? tmp_20_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_73 = _io_exe_rd_7_resp_T[21] ? tmp_21_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_74 = _io_exe_rd_7_resp_T[22] ? tmp_22_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_75 = _io_exe_rd_7_resp_T[23] ? tmp_23_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_76 = _io_exe_rd_7_resp_T[24] ? tmp_24_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_77 = _io_exe_rd_7_resp_T[25] ? tmp_25_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_78 = _io_exe_rd_7_resp_T[26] ? tmp_26_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_79 = _io_exe_rd_7_resp_T[27] ? tmp_27_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_80 = _io_exe_rd_7_resp_T[28] ? tmp_28_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_81 = _io_exe_rd_7_resp_T[29] ? tmp_29_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_82 = _io_exe_rd_7_resp_T[30] ? tmp_30_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_83 = _io_exe_rd_7_resp_T[31] ? tmp_31_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_84 = _io_exe_rd_7_resp_T[32] ? tmp_32_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_85 = _io_exe_rd_7_resp_T[33] ? tmp_33_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_86 = _io_exe_rd_7_resp_T[34] ? tmp_34_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_87 = _io_exe_rd_7_resp_T[35] ? tmp_35_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_88 = _io_exe_rd_7_resp_T[36] ? tmp_36_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_89 = _io_exe_rd_7_resp_T[37] ? tmp_37_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_90 = _io_exe_rd_7_resp_T[38] ? tmp_38_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_91 = _io_exe_rd_7_resp_T[39] ? tmp_39_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_92 = _io_exe_rd_7_resp_T[40] ? tmp_40_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_93 = _io_exe_rd_7_resp_T[41] ? tmp_41_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_94 = _io_exe_rd_7_resp_T[42] ? tmp_42_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_95 = _io_exe_rd_7_resp_T[43] ? tmp_43_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_96 = _io_exe_rd_7_resp_T[44] ? tmp_44_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_97 = _io_exe_rd_7_resp_T[45] ? tmp_45_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_98 = _io_exe_rd_7_resp_T[46] ? tmp_46_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_99 = _io_exe_rd_7_resp_T[47] ? tmp_47_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_100 = _io_exe_rd_7_resp_T[48] ? tmp_48_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_101 = _io_exe_rd_7_resp_T[49] ? tmp_49_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_102 = _io_exe_rd_7_resp_T[50] ? tmp_50_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_103 = _io_exe_rd_7_resp_T_52 | _io_exe_rd_7_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_104 = _io_exe_rd_7_resp_T_103 | _io_exe_rd_7_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_105 = _io_exe_rd_7_resp_T_104 | _io_exe_rd_7_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_106 = _io_exe_rd_7_resp_T_105 | _io_exe_rd_7_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_107 = _io_exe_rd_7_resp_T_106 | _io_exe_rd_7_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_108 = _io_exe_rd_7_resp_T_107 | _io_exe_rd_7_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_109 = _io_exe_rd_7_resp_T_108 | _io_exe_rd_7_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_110 = _io_exe_rd_7_resp_T_109 | _io_exe_rd_7_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_111 = _io_exe_rd_7_resp_T_110 | _io_exe_rd_7_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_112 = _io_exe_rd_7_resp_T_111 | _io_exe_rd_7_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_113 = _io_exe_rd_7_resp_T_112 | _io_exe_rd_7_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_114 = _io_exe_rd_7_resp_T_113 | _io_exe_rd_7_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_115 = _io_exe_rd_7_resp_T_114 | _io_exe_rd_7_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_116 = _io_exe_rd_7_resp_T_115 | _io_exe_rd_7_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_117 = _io_exe_rd_7_resp_T_116 | _io_exe_rd_7_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_118 = _io_exe_rd_7_resp_T_117 | _io_exe_rd_7_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_119 = _io_exe_rd_7_resp_T_118 | _io_exe_rd_7_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_120 = _io_exe_rd_7_resp_T_119 | _io_exe_rd_7_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_121 = _io_exe_rd_7_resp_T_120 | _io_exe_rd_7_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_122 = _io_exe_rd_7_resp_T_121 | _io_exe_rd_7_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_123 = _io_exe_rd_7_resp_T_122 | _io_exe_rd_7_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_124 = _io_exe_rd_7_resp_T_123 | _io_exe_rd_7_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_125 = _io_exe_rd_7_resp_T_124 | _io_exe_rd_7_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_126 = _io_exe_rd_7_resp_T_125 | _io_exe_rd_7_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_127 = _io_exe_rd_7_resp_T_126 | _io_exe_rd_7_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_128 = _io_exe_rd_7_resp_T_127 | _io_exe_rd_7_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_129 = _io_exe_rd_7_resp_T_128 | _io_exe_rd_7_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_130 = _io_exe_rd_7_resp_T_129 | _io_exe_rd_7_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_131 = _io_exe_rd_7_resp_T_130 | _io_exe_rd_7_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_132 = _io_exe_rd_7_resp_T_131 | _io_exe_rd_7_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_133 = _io_exe_rd_7_resp_T_132 | _io_exe_rd_7_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_134 = _io_exe_rd_7_resp_T_133 | _io_exe_rd_7_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_135 = _io_exe_rd_7_resp_T_134 | _io_exe_rd_7_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_136 = _io_exe_rd_7_resp_T_135 | _io_exe_rd_7_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_137 = _io_exe_rd_7_resp_T_136 | _io_exe_rd_7_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_138 = _io_exe_rd_7_resp_T_137 | _io_exe_rd_7_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_139 = _io_exe_rd_7_resp_T_138 | _io_exe_rd_7_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_140 = _io_exe_rd_7_resp_T_139 | _io_exe_rd_7_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_141 = _io_exe_rd_7_resp_T_140 | _io_exe_rd_7_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_142 = _io_exe_rd_7_resp_T_141 | _io_exe_rd_7_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_143 = _io_exe_rd_7_resp_T_142 | _io_exe_rd_7_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_144 = _io_exe_rd_7_resp_T_143 | _io_exe_rd_7_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_145 = _io_exe_rd_7_resp_T_144 | _io_exe_rd_7_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_146 = _io_exe_rd_7_resp_T_145 | _io_exe_rd_7_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_147 = _io_exe_rd_7_resp_T_146 | _io_exe_rd_7_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_148 = _io_exe_rd_7_resp_T_147 | _io_exe_rd_7_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_149 = _io_exe_rd_7_resp_T_148 | _io_exe_rd_7_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_150 = _io_exe_rd_7_resp_T_149 | _io_exe_rd_7_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_7_resp_T_151 = _io_exe_rd_7_resp_T_150 | _io_exe_rd_7_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_8 = io_exe_rd_8_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3665 = io_exe_rd_8_req_gidx[0] ? io_coef_in_mainch_drc_smooth_1 : io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h2 ? _GEN_3665 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_8 = io_exe_rd_8_req_iscoef ? tmp_8_out_out_out_8 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3669 = io_exe_rd_8_req_gidx[0] ? io_coef_in_subch_drc_smooth_1 : io_coef_in_subch_drc_smooth_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h2 ? _GEN_3669 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_8 = io_exe_rd_8_req_iscoef ? tmp_9_out_out_out_8 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3673 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3674 = 3'h2 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3673; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3675 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3674; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3676 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3675; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3676 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_8 = io_exe_rd_8_req_iscoef ? tmp_10_out_out_out_8 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_8 = io_exe_rd_8_req_iscoef ? tmp_10_out_out_out_8 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3687 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3688 = 3'h2 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3687; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3689 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3688; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3690 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3689; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3690 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_8 = io_exe_rd_8_req_iscoef ? tmp_12_out_out_out_8 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_8 = io_exe_rd_8_req_iscoef ? tmp_12_out_out_out_8 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3701 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3702 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_3701; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3703 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_3702; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3704 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_3703; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3704 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_34 = io_exe_rd_8_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_3707 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3708 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt__2 : _GEN_3707; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3709 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt__3 : _GEN_3708; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3709 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_14_out_out_out_17 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_8 = io_exe_rd_8_req_iscoef ? tmp_14_out_out_out_16 : tmp_14_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3714 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3715 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_3714; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3716 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_3715; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3717 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_3716; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3717 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3720 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3721 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_1_2 : _GEN_3720; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3722 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_1_3 : _GEN_3721; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3722 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_15_out_out_out_17 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_8 = io_exe_rd_8_req_iscoef ? tmp_15_out_out_out_16 : tmp_15_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3727 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3728 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_3727; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3729 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_3728; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3730 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_3729; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3730 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3733 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3734 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_2_2 : _GEN_3733; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3735 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_2_3 : _GEN_3734; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3735 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_16_out_out_out_17 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_8 = io_exe_rd_8_req_iscoef ? tmp_16_out_out_out_16 : tmp_16_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3740 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3741 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_3740; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3742 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_3741; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3743 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_3742; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3743 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3746 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3747 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_3_2 : _GEN_3746; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3748 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_3_3 : _GEN_3747; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3748 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_17_out_out_out_17 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_8 = io_exe_rd_8_req_iscoef ? tmp_17_out_out_out_16 : tmp_17_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3753 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3754 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_3753; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3755 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_3754; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3756 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_3755; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3756 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3759 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3760 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_4_2 : _GEN_3759; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3761 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_4_3 : _GEN_3760; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3761 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_18_out_out_out_17 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_8 = io_exe_rd_8_req_iscoef ? tmp_18_out_out_out_16 : tmp_18_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3766 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3767 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_3766; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3768 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_3767; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3769 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_3768; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3769 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3772 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3773 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_5_2 : _GEN_3772; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3774 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_5_3 : _GEN_3773; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3774 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_19_out_out_out_17 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_8 = io_exe_rd_8_req_iscoef ? tmp_19_out_out_out_16 : tmp_19_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3779 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3780 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_3779; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3781 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_3780; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3782 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_3781; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3782 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3785 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3786 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_6_2 : _GEN_3785; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3787 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_6_3 : _GEN_3786; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3787 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_20_out_out_out_17 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_8 = io_exe_rd_8_req_iscoef ? tmp_20_out_out_out_16 : tmp_20_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3792 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3793 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_3792; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3794 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_3793; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3795 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_3794; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3795 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3798 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3799 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_7_2 : _GEN_3798; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3800 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_7_3 : _GEN_3799; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3800 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_21_out_out_out_17 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_8 = io_exe_rd_8_req_iscoef ? tmp_21_out_out_out_16 : tmp_21_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3805 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3806 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_3805; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3807 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_3806; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3808 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_3807; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3808 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3811 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3812 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_8_2 : _GEN_3811; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3813 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_8_3 : _GEN_3812; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3813 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_22_out_out_out_17 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_8 = io_exe_rd_8_req_iscoef ? tmp_22_out_out_out_16 : tmp_22_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3818 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3819 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_3818; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3820 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_3819; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3821 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_3820; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3821 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3824 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3825 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_9_2 : _GEN_3824; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3826 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_9_3 : _GEN_3825; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3826 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_23_out_out_out_17 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_8 = io_exe_rd_8_req_iscoef ? tmp_23_out_out_out_16 : tmp_23_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3831 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3832 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_3831; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3833 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_3832; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3834 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_3833; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3834 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3837 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3838 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_10_2 : _GEN_3837; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3839 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_10_3 : _GEN_3838; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3839 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_24_out_out_out_17 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_8 = io_exe_rd_8_req_iscoef ? tmp_24_out_out_out_16 : tmp_24_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3844 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3845 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_3844; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3846 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_3845; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3847 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_3846; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3847 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3850 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3851 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_11_2 : _GEN_3850; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3852 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_11_3 : _GEN_3851; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3852 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_25_out_out_out_17 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_8 = io_exe_rd_8_req_iscoef ? tmp_25_out_out_out_16 : tmp_25_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3857 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3858 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_3857; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3859 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_3858; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3860 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_3859; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3860 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3863 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3864 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_12_2 : _GEN_3863; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3865 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_12_3 : _GEN_3864; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3865 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_26_out_out_out_17 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_8 = io_exe_rd_8_req_iscoef ? tmp_26_out_out_out_16 : tmp_26_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3870 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3871 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_3870; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3872 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_3871; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3873 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_3872; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3873 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3876 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3877 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_13_2 : _GEN_3876; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3878 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_13_3 : _GEN_3877; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3878 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_27_out_out_out_17 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_8 = io_exe_rd_8_req_iscoef ? tmp_27_out_out_out_16 : tmp_27_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3883 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3884 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_3883; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3885 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_3884; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3886 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_3885; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3886 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3889 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3890 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_14_2 : _GEN_3889; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3891 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_14_3 : _GEN_3890; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3891 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_28_out_out_out_17 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_8 = io_exe_rd_8_req_iscoef ? tmp_28_out_out_out_16 : tmp_28_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3896 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3897 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_3896; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3898 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_3897; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3899 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_3898; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3899 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3902 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3903 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_15_2 : _GEN_3902; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3904 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_15_3 : _GEN_3903; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3904 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_29_out_out_out_17 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_8 = io_exe_rd_8_req_iscoef ? tmp_29_out_out_out_16 : tmp_29_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3909 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3910 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_3909; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3911 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_3910; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3912 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_3911; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3912 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3915 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3916 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_16_2 : _GEN_3915; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3917 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_16_3 : _GEN_3916; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3917 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_30_out_out_out_17 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_8 = io_exe_rd_8_req_iscoef ? tmp_30_out_out_out_16 : tmp_30_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3922 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3923 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_3922; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3924 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_3923; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3925 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_3924; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3925 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3928 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3929 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_17_2 : _GEN_3928; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3930 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_17_3 : _GEN_3929; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3930 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_31_out_out_out_17 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_8 = io_exe_rd_8_req_iscoef ? tmp_31_out_out_out_16 : tmp_31_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3935 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3936 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_3935; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3937 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_3936; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3938 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_3937; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3938 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3941 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3942 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_18_2 : _GEN_3941; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3943 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_18_3 : _GEN_3942; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3943 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_32_out_out_out_17 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_8 = io_exe_rd_8_req_iscoef ? tmp_32_out_out_out_16 : tmp_32_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3948 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3949 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_3948; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3950 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_3949; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3951 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_3950; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3951 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3954 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3955 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_19_2 : _GEN_3954; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3956 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_19_3 : _GEN_3955; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3956 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_33_out_out_out_17 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_8 = io_exe_rd_8_req_iscoef ? tmp_33_out_out_out_16 : tmp_33_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3961 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3962 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_3961; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3963 = 3'h3 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_3962; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3964 = 3'h4 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_3963; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_16 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3964 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_3967 = 2'h1 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3968 = 2'h2 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_20_2 : _GEN_3967; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3969 = 2'h3 == _tmp_14_out_out_T_34[1:0] ? reg_type5_data_nxt_20_3 : _GEN_3968; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_17 = _tmp_14_out_out_T_34 < 3'h4 ? _GEN_3969 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_17 = io_exe_rd_8_req_isgroup ? tmp_34_out_out_out_17 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_8 = io_exe_rd_8_req_iscoef ? tmp_34_out_out_out_16 : tmp_34_out_out_17; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3974 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3975 = 3'h2 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3974; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3976 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3975; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3977 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3976; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3977 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_8 = io_exe_rd_8_req_iscoef ? tmp_35_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3981 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3982 = 3'h2 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3981; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3983 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3982; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3984 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3983; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3984 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_8 = io_exe_rd_8_req_iscoef ? tmp_36_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3988 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3989 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_3988; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3990 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3989; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3991 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3990; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3991 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_8 = io_exe_rd_8_req_iscoef ? tmp_37_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_3995 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3996 = 3'h2 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3995; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3997 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3996; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_3998 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_3997; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_3998 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_8 = io_exe_rd_8_req_iscoef ? tmp_38_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4002 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4003 = 3'h2 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4002; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4004 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4003; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4005 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4004; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_4005 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_8 = io_exe_rd_8_req_iscoef ? tmp_39_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4009 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4010 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_4009; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4011 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4010; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4012 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4011; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_4012 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_8 = io_exe_rd_8_req_iscoef ? tmp_40_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4016 = 3'h1 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4017 = 3'h2 == io_exe_rd_8_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_4016; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4018 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4017; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4019 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4018; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_4019 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_8 = io_exe_rd_8_req_iscoef ? tmp_41_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4023 = 3'h1 == io_exe_rd_8_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4024 = 3'h2 == io_exe_rd_8_req_gidx ? reg_type6_coef_7_2 : _GEN_4023; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4025 = 3'h3 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4024; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4026 = 3'h4 == io_exe_rd_8_req_gidx ? 32'h0 : _GEN_4025; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_8 = io_exe_rd_8_req_gidx < 3'h5 ? _GEN_4026 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_8 = io_exe_rd_8_req_iscoef ? tmp_42_out_out_out_8 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_8 = io_exe_rd_8_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_8 = io_exe_rd_8_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_8 = io_exe_rd_8_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_8 = io_exe_rd_8_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_8 = io_exe_rd_8_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_8 = io_exe_rd_8_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_8 = io_exe_rd_8_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_8 = io_exe_rd_8_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_8_resp_T = 64'h1 << io_exe_rd_8_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_8_resp_T_52 = _io_exe_rd_8_resp_T[0] ? tmp_0_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_53 = _io_exe_rd_8_resp_T[1] ? tmp_1_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_54 = _io_exe_rd_8_resp_T[2] ? tmp_2_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_55 = _io_exe_rd_8_resp_T[3] ? tmp_3_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_56 = _io_exe_rd_8_resp_T[4] ? tmp_4_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_57 = _io_exe_rd_8_resp_T[5] ? tmp_5_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_58 = _io_exe_rd_8_resp_T[6] ? tmp_6_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_59 = _io_exe_rd_8_resp_T[7] ? tmp_7_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_60 = _io_exe_rd_8_resp_T[8] ? tmp_8_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_61 = _io_exe_rd_8_resp_T[9] ? tmp_9_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_62 = _io_exe_rd_8_resp_T[10] ? tmp_10_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_63 = _io_exe_rd_8_resp_T[11] ? tmp_11_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_64 = _io_exe_rd_8_resp_T[12] ? tmp_12_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_65 = _io_exe_rd_8_resp_T[13] ? tmp_13_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_66 = _io_exe_rd_8_resp_T[14] ? tmp_14_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_67 = _io_exe_rd_8_resp_T[15] ? tmp_15_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_68 = _io_exe_rd_8_resp_T[16] ? tmp_16_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_69 = _io_exe_rd_8_resp_T[17] ? tmp_17_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_70 = _io_exe_rd_8_resp_T[18] ? tmp_18_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_71 = _io_exe_rd_8_resp_T[19] ? tmp_19_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_72 = _io_exe_rd_8_resp_T[20] ? tmp_20_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_73 = _io_exe_rd_8_resp_T[21] ? tmp_21_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_74 = _io_exe_rd_8_resp_T[22] ? tmp_22_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_75 = _io_exe_rd_8_resp_T[23] ? tmp_23_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_76 = _io_exe_rd_8_resp_T[24] ? tmp_24_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_77 = _io_exe_rd_8_resp_T[25] ? tmp_25_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_78 = _io_exe_rd_8_resp_T[26] ? tmp_26_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_79 = _io_exe_rd_8_resp_T[27] ? tmp_27_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_80 = _io_exe_rd_8_resp_T[28] ? tmp_28_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_81 = _io_exe_rd_8_resp_T[29] ? tmp_29_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_82 = _io_exe_rd_8_resp_T[30] ? tmp_30_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_83 = _io_exe_rd_8_resp_T[31] ? tmp_31_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_84 = _io_exe_rd_8_resp_T[32] ? tmp_32_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_85 = _io_exe_rd_8_resp_T[33] ? tmp_33_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_86 = _io_exe_rd_8_resp_T[34] ? tmp_34_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_87 = _io_exe_rd_8_resp_T[35] ? tmp_35_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_88 = _io_exe_rd_8_resp_T[36] ? tmp_36_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_89 = _io_exe_rd_8_resp_T[37] ? tmp_37_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_90 = _io_exe_rd_8_resp_T[38] ? tmp_38_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_91 = _io_exe_rd_8_resp_T[39] ? tmp_39_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_92 = _io_exe_rd_8_resp_T[40] ? tmp_40_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_93 = _io_exe_rd_8_resp_T[41] ? tmp_41_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_94 = _io_exe_rd_8_resp_T[42] ? tmp_42_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_95 = _io_exe_rd_8_resp_T[43] ? tmp_43_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_96 = _io_exe_rd_8_resp_T[44] ? tmp_44_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_97 = _io_exe_rd_8_resp_T[45] ? tmp_45_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_98 = _io_exe_rd_8_resp_T[46] ? tmp_46_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_99 = _io_exe_rd_8_resp_T[47] ? tmp_47_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_100 = _io_exe_rd_8_resp_T[48] ? tmp_48_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_101 = _io_exe_rd_8_resp_T[49] ? tmp_49_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_102 = _io_exe_rd_8_resp_T[50] ? tmp_50_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_103 = _io_exe_rd_8_resp_T_52 | _io_exe_rd_8_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_104 = _io_exe_rd_8_resp_T_103 | _io_exe_rd_8_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_105 = _io_exe_rd_8_resp_T_104 | _io_exe_rd_8_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_106 = _io_exe_rd_8_resp_T_105 | _io_exe_rd_8_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_107 = _io_exe_rd_8_resp_T_106 | _io_exe_rd_8_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_108 = _io_exe_rd_8_resp_T_107 | _io_exe_rd_8_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_109 = _io_exe_rd_8_resp_T_108 | _io_exe_rd_8_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_110 = _io_exe_rd_8_resp_T_109 | _io_exe_rd_8_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_111 = _io_exe_rd_8_resp_T_110 | _io_exe_rd_8_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_112 = _io_exe_rd_8_resp_T_111 | _io_exe_rd_8_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_113 = _io_exe_rd_8_resp_T_112 | _io_exe_rd_8_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_114 = _io_exe_rd_8_resp_T_113 | _io_exe_rd_8_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_115 = _io_exe_rd_8_resp_T_114 | _io_exe_rd_8_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_116 = _io_exe_rd_8_resp_T_115 | _io_exe_rd_8_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_117 = _io_exe_rd_8_resp_T_116 | _io_exe_rd_8_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_118 = _io_exe_rd_8_resp_T_117 | _io_exe_rd_8_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_119 = _io_exe_rd_8_resp_T_118 | _io_exe_rd_8_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_120 = _io_exe_rd_8_resp_T_119 | _io_exe_rd_8_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_121 = _io_exe_rd_8_resp_T_120 | _io_exe_rd_8_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_122 = _io_exe_rd_8_resp_T_121 | _io_exe_rd_8_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_123 = _io_exe_rd_8_resp_T_122 | _io_exe_rd_8_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_124 = _io_exe_rd_8_resp_T_123 | _io_exe_rd_8_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_125 = _io_exe_rd_8_resp_T_124 | _io_exe_rd_8_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_126 = _io_exe_rd_8_resp_T_125 | _io_exe_rd_8_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_127 = _io_exe_rd_8_resp_T_126 | _io_exe_rd_8_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_128 = _io_exe_rd_8_resp_T_127 | _io_exe_rd_8_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_129 = _io_exe_rd_8_resp_T_128 | _io_exe_rd_8_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_130 = _io_exe_rd_8_resp_T_129 | _io_exe_rd_8_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_131 = _io_exe_rd_8_resp_T_130 | _io_exe_rd_8_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_132 = _io_exe_rd_8_resp_T_131 | _io_exe_rd_8_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_133 = _io_exe_rd_8_resp_T_132 | _io_exe_rd_8_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_134 = _io_exe_rd_8_resp_T_133 | _io_exe_rd_8_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_135 = _io_exe_rd_8_resp_T_134 | _io_exe_rd_8_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_136 = _io_exe_rd_8_resp_T_135 | _io_exe_rd_8_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_137 = _io_exe_rd_8_resp_T_136 | _io_exe_rd_8_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_138 = _io_exe_rd_8_resp_T_137 | _io_exe_rd_8_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_139 = _io_exe_rd_8_resp_T_138 | _io_exe_rd_8_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_140 = _io_exe_rd_8_resp_T_139 | _io_exe_rd_8_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_141 = _io_exe_rd_8_resp_T_140 | _io_exe_rd_8_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_142 = _io_exe_rd_8_resp_T_141 | _io_exe_rd_8_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_143 = _io_exe_rd_8_resp_T_142 | _io_exe_rd_8_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_144 = _io_exe_rd_8_resp_T_143 | _io_exe_rd_8_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_145 = _io_exe_rd_8_resp_T_144 | _io_exe_rd_8_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_146 = _io_exe_rd_8_resp_T_145 | _io_exe_rd_8_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_147 = _io_exe_rd_8_resp_T_146 | _io_exe_rd_8_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_148 = _io_exe_rd_8_resp_T_147 | _io_exe_rd_8_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_149 = _io_exe_rd_8_resp_T_148 | _io_exe_rd_8_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_150 = _io_exe_rd_8_resp_T_149 | _io_exe_rd_8_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_8_resp_T_151 = _io_exe_rd_8_resp_T_150 | _io_exe_rd_8_resp_T_101; // @[Mux.scala 27:72]
  wire [31:0] tmp_0_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type1_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_1_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type1_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_2_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type1_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_3_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type1_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_4_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type2_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_5_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type2_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_6_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type2_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_7_out_9 = io_exe_rd_9_req_iscoef ? 32'h0 : reg_type2_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_8_out_coef_out_9_0 = io_exe_rd_9_req_sel ? io_coef_in_mainch_drc_smooth_2 :
    io_coef_in_mainch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_8_out_coef_out_9_1 = io_exe_rd_9_req_sel ? io_coef_in_mainch_drc_smooth_3 :
    io_coef_in_mainch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_4046 = io_exe_rd_9_req_gidx[0] ? tmp_8_out_coef_out_9_1 : tmp_8_out_coef_out_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_8_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h2 ? _GEN_4046 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_8_out_9 = io_exe_rd_9_req_iscoef ? tmp_8_out_out_out_9 : reg_type3_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_9_out_coef_out_9_0 = io_exe_rd_9_req_sel ? io_coef_in_subch_drc_smooth_2 :
    io_coef_in_subch_drc_smooth_0; // @[regfile.scala 88:29]
  wire [31:0] tmp_9_out_coef_out_9_1 = io_exe_rd_9_req_sel ? io_coef_in_subch_drc_smooth_3 :
    io_coef_in_subch_drc_smooth_1; // @[regfile.scala 89:29]
  wire [31:0] _GEN_4050 = io_exe_rd_9_req_gidx[0] ? tmp_9_out_coef_out_9_1 : tmp_9_out_coef_out_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_9_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h2 ? _GEN_4050 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_9_out_9 = io_exe_rd_9_req_iscoef ? tmp_9_out_out_out_9 : reg_type3_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4054 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_drc_pow_1 : io_coef_in_mainch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4055 = 3'h2 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4054; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4056 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4055; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4057 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4056; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_10_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4057 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_10_out_9 = io_exe_rd_9_req_iscoef ? tmp_10_out_out_out_9 : reg_type4_data_nxt_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_11_out_9 = io_exe_rd_9_req_iscoef ? tmp_10_out_out_out_9 : reg_type4_data_nxt_1_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4068 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_subch_drc_pow_1 : io_coef_in_subch_drc_pow_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4069 = 3'h2 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4068; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4070 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4069; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4071 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4070; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_12_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4071 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_12_out_9 = io_exe_rd_9_req_iscoef ? tmp_12_out_out_out_9 : reg_type4_data_nxt_2_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_13_out_9 = io_exe_rd_9_req_iscoef ? tmp_12_out_out_out_9 : reg_type4_data_nxt_3_0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4082 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_1 :
    io_coef_in_mainch_ch0_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4083 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_2 : _GEN_4082; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4084 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_3 : _GEN_4083; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4085 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_0_4 : _GEN_4084; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4085 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [2:0] _tmp_14_out_out_T_38 = io_exe_rd_9_req_gidx - 3'h1; // @[regfile.scala 71:37]
  wire [31:0] _GEN_4088 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt__1 : reg_type5_data_nxt__0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4089 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt__2 : _GEN_4088; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4090 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt__3 : _GEN_4089; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4090 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_14_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_14_out_out_out_19 : reg_type5_data_nxt__2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_14_out_9 = io_exe_rd_9_req_iscoef ? tmp_14_out_out_out_18 : tmp_14_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4095 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_1 :
    io_coef_in_mainch_ch0_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4096 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_2 : _GEN_4095; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4097 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_3 : _GEN_4096; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4098 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_1_4 : _GEN_4097; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4098 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4101 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_1_1 : reg_type5_data_nxt_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4102 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_1_2 : _GEN_4101; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4103 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_1_3 : _GEN_4102; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4103 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_15_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_15_out_out_out_19 : reg_type5_data_nxt_1_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_15_out_9 = io_exe_rd_9_req_iscoef ? tmp_15_out_out_out_18 : tmp_15_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4108 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_1 :
    io_coef_in_mainch_ch0_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4109 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_2 : _GEN_4108; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4110 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_3 : _GEN_4109; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4111 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_2_4 : _GEN_4110; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4111 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4114 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_2_1 : reg_type5_data_nxt_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4115 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_2_2 : _GEN_4114; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4116 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_2_3 : _GEN_4115; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4116 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_16_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_16_out_out_out_19 : reg_type5_data_nxt_2_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_16_out_9 = io_exe_rd_9_req_iscoef ? tmp_16_out_out_out_18 : tmp_16_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4121 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_1 :
    io_coef_in_mainch_ch0_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4122 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_2 : _GEN_4121; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4123 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_3 : _GEN_4122; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4124 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_3_4 : _GEN_4123; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4124 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4127 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_3_1 : reg_type5_data_nxt_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4128 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_3_2 : _GEN_4127; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4129 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_3_3 : _GEN_4128; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4129 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_17_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_17_out_out_out_19 : reg_type5_data_nxt_3_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_17_out_9 = io_exe_rd_9_req_iscoef ? tmp_17_out_out_out_18 : tmp_17_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4134 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_1 :
    io_coef_in_mainch_ch0_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4135 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_2 : _GEN_4134; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4136 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_3 : _GEN_4135; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4137 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_4_4 : _GEN_4136; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4137 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4140 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_4_1 : reg_type5_data_nxt_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4141 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_4_2 : _GEN_4140; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4142 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_4_3 : _GEN_4141; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4142 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_18_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_18_out_out_out_19 : reg_type5_data_nxt_4_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_18_out_9 = io_exe_rd_9_req_iscoef ? tmp_18_out_out_out_18 : tmp_18_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4147 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_1 :
    io_coef_in_mainch_ch0_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4148 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_2 : _GEN_4147; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4149 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_3 : _GEN_4148; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4150 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_5_4 : _GEN_4149; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4150 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4153 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_5_1 : reg_type5_data_nxt_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4154 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_5_2 : _GEN_4153; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4155 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_5_3 : _GEN_4154; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4155 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_19_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_19_out_out_out_19 : reg_type5_data_nxt_5_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_19_out_9 = io_exe_rd_9_req_iscoef ? tmp_19_out_out_out_18 : tmp_19_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4160 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_1 :
    io_coef_in_mainch_ch0_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4161 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_2 : _GEN_4160; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4162 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_3 : _GEN_4161; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4163 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_6_4 : _GEN_4162; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4163 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4166 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_6_1 : reg_type5_data_nxt_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4167 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_6_2 : _GEN_4166; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4168 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_6_3 : _GEN_4167; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4168 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_20_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_20_out_out_out_19 : reg_type5_data_nxt_6_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_20_out_9 = io_exe_rd_9_req_iscoef ? tmp_20_out_out_out_18 : tmp_20_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4173 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_1 :
    io_coef_in_mainch_ch0_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4174 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_2 : _GEN_4173; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4175 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_3 : _GEN_4174; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4176 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_7_4 : _GEN_4175; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4176 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4179 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_7_1 : reg_type5_data_nxt_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4180 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_7_2 : _GEN_4179; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4181 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_7_3 : _GEN_4180; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4181 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_21_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_21_out_out_out_19 : reg_type5_data_nxt_7_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_21_out_9 = io_exe_rd_9_req_iscoef ? tmp_21_out_out_out_18 : tmp_21_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4186 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_1 :
    io_coef_in_mainch_ch0_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4187 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_2 : _GEN_4186; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4188 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_3 : _GEN_4187; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4189 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_bqcoef_8_4 : _GEN_4188; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4189 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4192 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_8_1 : reg_type5_data_nxt_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4193 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_8_2 : _GEN_4192; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4194 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_8_3 : _GEN_4193; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4194 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_22_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_22_out_out_out_19 : reg_type5_data_nxt_8_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_22_out_9 = io_exe_rd_9_req_iscoef ? tmp_22_out_out_out_18 : tmp_22_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4199 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_1 :
    io_coef_in_mainch_ch1_bqcoef_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4200 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_2 : _GEN_4199; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4201 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_3 : _GEN_4200; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4202 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_0_4 : _GEN_4201; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4202 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4205 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_9_1 : reg_type5_data_nxt_9_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4206 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_9_2 : _GEN_4205; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4207 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_9_3 : _GEN_4206; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4207 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_23_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_23_out_out_out_19 : reg_type5_data_nxt_9_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_23_out_9 = io_exe_rd_9_req_iscoef ? tmp_23_out_out_out_18 : tmp_23_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4212 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_1 :
    io_coef_in_mainch_ch1_bqcoef_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4213 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_2 : _GEN_4212; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4214 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_3 : _GEN_4213; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4215 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_1_4 : _GEN_4214; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4215 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4218 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_10_1 : reg_type5_data_nxt_10_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4219 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_10_2 : _GEN_4218; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4220 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_10_3 : _GEN_4219; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4220 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_24_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_24_out_out_out_19 : reg_type5_data_nxt_10_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_24_out_9 = io_exe_rd_9_req_iscoef ? tmp_24_out_out_out_18 : tmp_24_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4225 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_1 :
    io_coef_in_mainch_ch1_bqcoef_2_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4226 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_2 : _GEN_4225; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4227 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_3 : _GEN_4226; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4228 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_2_4 : _GEN_4227; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4228 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4231 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_11_1 : reg_type5_data_nxt_11_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4232 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_11_2 : _GEN_4231; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4233 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_11_3 : _GEN_4232; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4233 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_25_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_25_out_out_out_19 : reg_type5_data_nxt_11_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_25_out_9 = io_exe_rd_9_req_iscoef ? tmp_25_out_out_out_18 : tmp_25_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4238 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_1 :
    io_coef_in_mainch_ch1_bqcoef_3_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4239 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_2 : _GEN_4238; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4240 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_3 : _GEN_4239; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4241 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_3_4 : _GEN_4240; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4241 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4244 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_12_1 : reg_type5_data_nxt_12_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4245 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_12_2 : _GEN_4244; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4246 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_12_3 : _GEN_4245; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4246 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_26_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_26_out_out_out_19 : reg_type5_data_nxt_12_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_26_out_9 = io_exe_rd_9_req_iscoef ? tmp_26_out_out_out_18 : tmp_26_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4251 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_1 :
    io_coef_in_mainch_ch1_bqcoef_4_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4252 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_2 : _GEN_4251; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4253 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_3 : _GEN_4252; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4254 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_4_4 : _GEN_4253; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4254 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4257 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_13_1 : reg_type5_data_nxt_13_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4258 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_13_2 : _GEN_4257; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4259 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_13_3 : _GEN_4258; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4259 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_27_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_27_out_out_out_19 : reg_type5_data_nxt_13_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_27_out_9 = io_exe_rd_9_req_iscoef ? tmp_27_out_out_out_18 : tmp_27_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4264 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_1 :
    io_coef_in_mainch_ch1_bqcoef_5_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4265 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_2 : _GEN_4264; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4266 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_3 : _GEN_4265; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4267 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_5_4 : _GEN_4266; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4267 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4270 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_14_1 : reg_type5_data_nxt_14_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4271 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_14_2 : _GEN_4270; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4272 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_14_3 : _GEN_4271; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4272 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_28_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_28_out_out_out_19 : reg_type5_data_nxt_14_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_28_out_9 = io_exe_rd_9_req_iscoef ? tmp_28_out_out_out_18 : tmp_28_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4277 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_1 :
    io_coef_in_mainch_ch1_bqcoef_6_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4278 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_2 : _GEN_4277; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4279 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_3 : _GEN_4278; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4280 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_6_4 : _GEN_4279; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4280 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4283 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_15_1 : reg_type5_data_nxt_15_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4284 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_15_2 : _GEN_4283; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4285 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_15_3 : _GEN_4284; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4285 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_29_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_29_out_out_out_19 : reg_type5_data_nxt_15_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_29_out_9 = io_exe_rd_9_req_iscoef ? tmp_29_out_out_out_18 : tmp_29_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4290 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_1 :
    io_coef_in_mainch_ch1_bqcoef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4291 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_2 : _GEN_4290; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4292 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_3 : _GEN_4291; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4293 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_7_4 : _GEN_4292; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4293 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4296 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_16_1 : reg_type5_data_nxt_16_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4297 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_16_2 : _GEN_4296; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4298 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_16_3 : _GEN_4297; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4298 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_30_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_30_out_out_out_19 : reg_type5_data_nxt_16_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_30_out_9 = io_exe_rd_9_req_iscoef ? tmp_30_out_out_out_18 : tmp_30_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4303 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_1 :
    io_coef_in_mainch_ch1_bqcoef_8_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4304 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_2 : _GEN_4303; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4305 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_3 : _GEN_4304; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4306 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_bqcoef_8_4 : _GEN_4305; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4306 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4309 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_17_1 : reg_type5_data_nxt_17_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4310 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_17_2 : _GEN_4309; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4311 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_17_3 : _GEN_4310; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4311 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_31_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_31_out_out_out_19 : reg_type5_data_nxt_17_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_31_out_9 = io_exe_rd_9_req_iscoef ? tmp_31_out_out_out_18 : tmp_31_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4316 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch2bq_0_1 : io_coef_in_subch_ch2bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4317 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch2bq_0_2 : _GEN_4316; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4318 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch2bq_0_3 : _GEN_4317; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4319 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch2bq_0_4 : _GEN_4318; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4319 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4322 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_18_1 : reg_type5_data_nxt_18_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4323 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_18_2 : _GEN_4322; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4324 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_18_3 : _GEN_4323; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4324 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_32_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_32_out_out_out_19 : reg_type5_data_nxt_18_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_32_out_9 = io_exe_rd_9_req_iscoef ? tmp_32_out_out_out_18 : tmp_32_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4329 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_0_1 : io_coef_in_subch_ch3bq_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4330 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_0_2 : _GEN_4329; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4331 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_0_3 : _GEN_4330; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4332 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_0_4 : _GEN_4331; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4332 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4335 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_19_1 : reg_type5_data_nxt_19_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4336 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_19_2 : _GEN_4335; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4337 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_19_3 : _GEN_4336; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4337 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_33_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_33_out_out_out_19 : reg_type5_data_nxt_19_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_33_out_9 = io_exe_rd_9_req_iscoef ? tmp_33_out_out_out_18 : tmp_33_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4342 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_1_1 : io_coef_in_subch_ch3bq_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4343 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_1_2 : _GEN_4342; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4344 = 3'h3 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_1_3 : _GEN_4343; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4345 = 3'h4 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch3bq_1_4 : _GEN_4344; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_18 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4345 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] _GEN_4348 = 2'h1 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_20_1 : reg_type5_data_nxt_20_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4349 = 2'h2 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_20_2 : _GEN_4348; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4350 = 2'h3 == _tmp_14_out_out_T_38[1:0] ? reg_type5_data_nxt_20_3 : _GEN_4349; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_out_19 = _tmp_14_out_out_T_38 < 3'h4 ? _GEN_4350 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_34_out_out_19 = io_exe_rd_9_req_isgroup ? tmp_34_out_out_out_19 : reg_type5_data_nxt_20_2; // @[regfile.scala 70:27 regfile.scala 71:15 regfile.scala 73:15]
  wire [31:0] tmp_34_out_9 = io_exe_rd_9_req_iscoef ? tmp_34_out_out_out_18 : tmp_34_out_out_19; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4355 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_inputmix_0_1 :
    io_coef_in_mainch_ch0_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4356 = 3'h2 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4355; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4357 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4356; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4358 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4357; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_35_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4358 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_35_out_9 = io_exe_rd_9_req_iscoef ? tmp_35_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4362 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_inputmix_1_1 :
    io_coef_in_mainch_ch0_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4363 = 3'h2 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4362; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4364 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4363; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4365 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4364; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_36_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4365 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_36_out_9 = io_exe_rd_9_req_iscoef ? tmp_36_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4369 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_outputmix_1 :
    io_coef_in_mainch_ch0_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4370 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch0_outputmix_2 : _GEN_4369; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4371 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4370; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4372 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4371; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_37_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4372 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_37_out_9 = io_exe_rd_9_req_iscoef ? tmp_37_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4376 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_inputmix_0_1 :
    io_coef_in_mainch_ch1_inputmix_0_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4377 = 3'h2 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4376; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4378 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4377; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4379 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4378; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_38_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4379 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_38_out_9 = io_exe_rd_9_req_iscoef ? tmp_38_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4383 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_inputmix_1_1 :
    io_coef_in_mainch_ch1_inputmix_1_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4384 = 3'h2 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4383; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4385 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4384; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4386 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4385; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_39_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4386 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_39_out_9 = io_exe_rd_9_req_iscoef ? tmp_39_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4390 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_outputmix_1 :
    io_coef_in_mainch_ch1_outputmix_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4391 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_mainch_ch1_outputmix_2 : _GEN_4390; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4392 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4391; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4393 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4392; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_40_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4393 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_40_out_9 = io_exe_rd_9_req_iscoef ? tmp_40_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4397 = 3'h1 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch2mix_1 : io_coef_in_subch_ch2mix_2; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4398 = 3'h2 == io_exe_rd_9_req_gidx ? io_coef_in_subch_ch2mix_0 : _GEN_4397; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4399 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4398; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4400 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4399; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_41_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4400 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_41_out_9 = io_exe_rd_9_req_iscoef ? tmp_41_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] _GEN_4404 = 3'h1 == io_exe_rd_9_req_gidx ? reg_type6_coef_7_1 : reg_type6_coef_7_0; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4405 = 3'h2 == io_exe_rd_9_req_gidx ? reg_type6_coef_7_2 : _GEN_4404; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4406 = 3'h3 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4405; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] _GEN_4407 = 3'h4 == io_exe_rd_9_req_gidx ? 32'h0 : _GEN_4406; // @[regfile.scala 33:11 regfile.scala 33:11]
  wire [31:0] tmp_42_out_out_out_9 = io_exe_rd_9_req_gidx < 3'h5 ? _GEN_4407 : 32'h0; // @[regfile.scala 32:29 regfile.scala 33:11]
  wire [31:0] tmp_42_out_9 = io_exe_rd_9_req_iscoef ? tmp_42_out_out_out_9 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_43_out_9 = io_exe_rd_9_req_iscoef ? io_coef_in_mainch_ch0_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_44_out_9 = io_exe_rd_9_req_iscoef ? io_coef_in_mainch_ch1_vol : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_45_out_9 = io_exe_rd_9_req_iscoef ? reg_type7_coef_2_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_46_out_9 = io_exe_rd_9_req_iscoef ? reg_type7_coef_3_0 : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_47_out_9 = io_exe_rd_9_req_iscoef ? io_coef_in_mainch_ch0_prescale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_48_out_9 = io_exe_rd_9_req_iscoef ? io_coef_in_mainch_ch0_postscale : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_49_out_9 = io_exe_rd_9_req_iscoef ? io_coef_in_mainch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [31:0] tmp_50_out_9 = io_exe_rd_9_req_iscoef ? io_coef_in_subch_drc_ratio : 32'h0; // @[regfile.scala 103:22 regfile.scala 104:11 regfile.scala 106:11]
  wire [63:0] _io_exe_rd_9_resp_T = 64'h1 << io_exe_rd_9_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_9_resp_T_52 = _io_exe_rd_9_resp_T[0] ? tmp_0_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_53 = _io_exe_rd_9_resp_T[1] ? tmp_1_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_54 = _io_exe_rd_9_resp_T[2] ? tmp_2_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_55 = _io_exe_rd_9_resp_T[3] ? tmp_3_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_56 = _io_exe_rd_9_resp_T[4] ? tmp_4_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_57 = _io_exe_rd_9_resp_T[5] ? tmp_5_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_58 = _io_exe_rd_9_resp_T[6] ? tmp_6_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_59 = _io_exe_rd_9_resp_T[7] ? tmp_7_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_60 = _io_exe_rd_9_resp_T[8] ? tmp_8_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_61 = _io_exe_rd_9_resp_T[9] ? tmp_9_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_62 = _io_exe_rd_9_resp_T[10] ? tmp_10_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_63 = _io_exe_rd_9_resp_T[11] ? tmp_11_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_64 = _io_exe_rd_9_resp_T[12] ? tmp_12_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_65 = _io_exe_rd_9_resp_T[13] ? tmp_13_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_66 = _io_exe_rd_9_resp_T[14] ? tmp_14_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_67 = _io_exe_rd_9_resp_T[15] ? tmp_15_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_68 = _io_exe_rd_9_resp_T[16] ? tmp_16_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_69 = _io_exe_rd_9_resp_T[17] ? tmp_17_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_70 = _io_exe_rd_9_resp_T[18] ? tmp_18_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_71 = _io_exe_rd_9_resp_T[19] ? tmp_19_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_72 = _io_exe_rd_9_resp_T[20] ? tmp_20_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_73 = _io_exe_rd_9_resp_T[21] ? tmp_21_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_74 = _io_exe_rd_9_resp_T[22] ? tmp_22_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_75 = _io_exe_rd_9_resp_T[23] ? tmp_23_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_76 = _io_exe_rd_9_resp_T[24] ? tmp_24_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_77 = _io_exe_rd_9_resp_T[25] ? tmp_25_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_78 = _io_exe_rd_9_resp_T[26] ? tmp_26_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_79 = _io_exe_rd_9_resp_T[27] ? tmp_27_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_80 = _io_exe_rd_9_resp_T[28] ? tmp_28_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_81 = _io_exe_rd_9_resp_T[29] ? tmp_29_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_82 = _io_exe_rd_9_resp_T[30] ? tmp_30_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_83 = _io_exe_rd_9_resp_T[31] ? tmp_31_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_84 = _io_exe_rd_9_resp_T[32] ? tmp_32_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_85 = _io_exe_rd_9_resp_T[33] ? tmp_33_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_86 = _io_exe_rd_9_resp_T[34] ? tmp_34_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_87 = _io_exe_rd_9_resp_T[35] ? tmp_35_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_88 = _io_exe_rd_9_resp_T[36] ? tmp_36_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_89 = _io_exe_rd_9_resp_T[37] ? tmp_37_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_90 = _io_exe_rd_9_resp_T[38] ? tmp_38_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_91 = _io_exe_rd_9_resp_T[39] ? tmp_39_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_92 = _io_exe_rd_9_resp_T[40] ? tmp_40_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_93 = _io_exe_rd_9_resp_T[41] ? tmp_41_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_94 = _io_exe_rd_9_resp_T[42] ? tmp_42_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_95 = _io_exe_rd_9_resp_T[43] ? tmp_43_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_96 = _io_exe_rd_9_resp_T[44] ? tmp_44_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_97 = _io_exe_rd_9_resp_T[45] ? tmp_45_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_98 = _io_exe_rd_9_resp_T[46] ? tmp_46_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_99 = _io_exe_rd_9_resp_T[47] ? tmp_47_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_100 = _io_exe_rd_9_resp_T[48] ? tmp_48_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_101 = _io_exe_rd_9_resp_T[49] ? tmp_49_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_102 = _io_exe_rd_9_resp_T[50] ? tmp_50_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_103 = _io_exe_rd_9_resp_T_52 | _io_exe_rd_9_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_104 = _io_exe_rd_9_resp_T_103 | _io_exe_rd_9_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_105 = _io_exe_rd_9_resp_T_104 | _io_exe_rd_9_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_106 = _io_exe_rd_9_resp_T_105 | _io_exe_rd_9_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_107 = _io_exe_rd_9_resp_T_106 | _io_exe_rd_9_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_108 = _io_exe_rd_9_resp_T_107 | _io_exe_rd_9_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_109 = _io_exe_rd_9_resp_T_108 | _io_exe_rd_9_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_110 = _io_exe_rd_9_resp_T_109 | _io_exe_rd_9_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_111 = _io_exe_rd_9_resp_T_110 | _io_exe_rd_9_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_112 = _io_exe_rd_9_resp_T_111 | _io_exe_rd_9_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_113 = _io_exe_rd_9_resp_T_112 | _io_exe_rd_9_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_114 = _io_exe_rd_9_resp_T_113 | _io_exe_rd_9_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_115 = _io_exe_rd_9_resp_T_114 | _io_exe_rd_9_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_116 = _io_exe_rd_9_resp_T_115 | _io_exe_rd_9_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_117 = _io_exe_rd_9_resp_T_116 | _io_exe_rd_9_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_118 = _io_exe_rd_9_resp_T_117 | _io_exe_rd_9_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_119 = _io_exe_rd_9_resp_T_118 | _io_exe_rd_9_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_120 = _io_exe_rd_9_resp_T_119 | _io_exe_rd_9_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_121 = _io_exe_rd_9_resp_T_120 | _io_exe_rd_9_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_122 = _io_exe_rd_9_resp_T_121 | _io_exe_rd_9_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_123 = _io_exe_rd_9_resp_T_122 | _io_exe_rd_9_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_124 = _io_exe_rd_9_resp_T_123 | _io_exe_rd_9_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_125 = _io_exe_rd_9_resp_T_124 | _io_exe_rd_9_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_126 = _io_exe_rd_9_resp_T_125 | _io_exe_rd_9_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_127 = _io_exe_rd_9_resp_T_126 | _io_exe_rd_9_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_128 = _io_exe_rd_9_resp_T_127 | _io_exe_rd_9_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_129 = _io_exe_rd_9_resp_T_128 | _io_exe_rd_9_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_130 = _io_exe_rd_9_resp_T_129 | _io_exe_rd_9_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_131 = _io_exe_rd_9_resp_T_130 | _io_exe_rd_9_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_132 = _io_exe_rd_9_resp_T_131 | _io_exe_rd_9_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_133 = _io_exe_rd_9_resp_T_132 | _io_exe_rd_9_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_134 = _io_exe_rd_9_resp_T_133 | _io_exe_rd_9_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_135 = _io_exe_rd_9_resp_T_134 | _io_exe_rd_9_resp_T_85; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_136 = _io_exe_rd_9_resp_T_135 | _io_exe_rd_9_resp_T_86; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_137 = _io_exe_rd_9_resp_T_136 | _io_exe_rd_9_resp_T_87; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_138 = _io_exe_rd_9_resp_T_137 | _io_exe_rd_9_resp_T_88; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_139 = _io_exe_rd_9_resp_T_138 | _io_exe_rd_9_resp_T_89; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_140 = _io_exe_rd_9_resp_T_139 | _io_exe_rd_9_resp_T_90; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_141 = _io_exe_rd_9_resp_T_140 | _io_exe_rd_9_resp_T_91; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_142 = _io_exe_rd_9_resp_T_141 | _io_exe_rd_9_resp_T_92; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_143 = _io_exe_rd_9_resp_T_142 | _io_exe_rd_9_resp_T_93; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_144 = _io_exe_rd_9_resp_T_143 | _io_exe_rd_9_resp_T_94; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_145 = _io_exe_rd_9_resp_T_144 | _io_exe_rd_9_resp_T_95; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_146 = _io_exe_rd_9_resp_T_145 | _io_exe_rd_9_resp_T_96; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_147 = _io_exe_rd_9_resp_T_146 | _io_exe_rd_9_resp_T_97; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_148 = _io_exe_rd_9_resp_T_147 | _io_exe_rd_9_resp_T_98; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_149 = _io_exe_rd_9_resp_T_148 | _io_exe_rd_9_resp_T_99; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_150 = _io_exe_rd_9_resp_T_149 | _io_exe_rd_9_resp_T_100; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_9_resp_T_151 = _io_exe_rd_9_resp_T_150 | _io_exe_rd_9_resp_T_101; // @[Mux.scala 27:72]
  wire [63:0] _io_exe_rd_10_resp_T = 64'h1 << io_exe_rd_10_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_10_resp_T_52 = _io_exe_rd_10_resp_T[0] ? reg_type1_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_53 = _io_exe_rd_10_resp_T[1] ? reg_type1_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_54 = _io_exe_rd_10_resp_T[2] ? reg_type1_data_nxt_2_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_55 = _io_exe_rd_10_resp_T[3] ? reg_type1_data_nxt_3_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_56 = _io_exe_rd_10_resp_T[4] ? reg_type2_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_57 = _io_exe_rd_10_resp_T[5] ? reg_type2_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_58 = _io_exe_rd_10_resp_T[6] ? reg_type2_data_nxt_2_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_59 = _io_exe_rd_10_resp_T[7] ? reg_type2_data_nxt_3_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_60 = _io_exe_rd_10_resp_T[8] ? reg_type3_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_61 = _io_exe_rd_10_resp_T[9] ? reg_type3_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_62 = _io_exe_rd_10_resp_T[10] ? reg_type4_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_63 = _io_exe_rd_10_resp_T[11] ? reg_type4_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_64 = _io_exe_rd_10_resp_T[12] ? reg_type4_data_nxt_2_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_65 = _io_exe_rd_10_resp_T[13] ? reg_type4_data_nxt_3_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_66 = _io_exe_rd_10_resp_T[14] ? reg_type5_data_nxt__2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_67 = _io_exe_rd_10_resp_T[15] ? reg_type5_data_nxt_1_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_68 = _io_exe_rd_10_resp_T[16] ? reg_type5_data_nxt_2_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_69 = _io_exe_rd_10_resp_T[17] ? reg_type5_data_nxt_3_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_70 = _io_exe_rd_10_resp_T[18] ? reg_type5_data_nxt_4_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_71 = _io_exe_rd_10_resp_T[19] ? reg_type5_data_nxt_5_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_72 = _io_exe_rd_10_resp_T[20] ? reg_type5_data_nxt_6_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_73 = _io_exe_rd_10_resp_T[21] ? reg_type5_data_nxt_7_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_74 = _io_exe_rd_10_resp_T[22] ? reg_type5_data_nxt_8_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_75 = _io_exe_rd_10_resp_T[23] ? reg_type5_data_nxt_9_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_76 = _io_exe_rd_10_resp_T[24] ? reg_type5_data_nxt_10_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_77 = _io_exe_rd_10_resp_T[25] ? reg_type5_data_nxt_11_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_78 = _io_exe_rd_10_resp_T[26] ? reg_type5_data_nxt_12_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_79 = _io_exe_rd_10_resp_T[27] ? reg_type5_data_nxt_13_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_80 = _io_exe_rd_10_resp_T[28] ? reg_type5_data_nxt_14_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_81 = _io_exe_rd_10_resp_T[29] ? reg_type5_data_nxt_15_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_82 = _io_exe_rd_10_resp_T[30] ? reg_type5_data_nxt_16_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_83 = _io_exe_rd_10_resp_T[31] ? reg_type5_data_nxt_17_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_84 = _io_exe_rd_10_resp_T[32] ? reg_type5_data_nxt_18_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_85 = _io_exe_rd_10_resp_T[33] ? reg_type5_data_nxt_19_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_86 = _io_exe_rd_10_resp_T[34] ? reg_type5_data_nxt_20_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_103 = _io_exe_rd_10_resp_T_52 | _io_exe_rd_10_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_104 = _io_exe_rd_10_resp_T_103 | _io_exe_rd_10_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_105 = _io_exe_rd_10_resp_T_104 | _io_exe_rd_10_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_106 = _io_exe_rd_10_resp_T_105 | _io_exe_rd_10_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_107 = _io_exe_rd_10_resp_T_106 | _io_exe_rd_10_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_108 = _io_exe_rd_10_resp_T_107 | _io_exe_rd_10_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_109 = _io_exe_rd_10_resp_T_108 | _io_exe_rd_10_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_110 = _io_exe_rd_10_resp_T_109 | _io_exe_rd_10_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_111 = _io_exe_rd_10_resp_T_110 | _io_exe_rd_10_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_112 = _io_exe_rd_10_resp_T_111 | _io_exe_rd_10_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_113 = _io_exe_rd_10_resp_T_112 | _io_exe_rd_10_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_114 = _io_exe_rd_10_resp_T_113 | _io_exe_rd_10_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_115 = _io_exe_rd_10_resp_T_114 | _io_exe_rd_10_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_116 = _io_exe_rd_10_resp_T_115 | _io_exe_rd_10_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_117 = _io_exe_rd_10_resp_T_116 | _io_exe_rd_10_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_118 = _io_exe_rd_10_resp_T_117 | _io_exe_rd_10_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_119 = _io_exe_rd_10_resp_T_118 | _io_exe_rd_10_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_120 = _io_exe_rd_10_resp_T_119 | _io_exe_rd_10_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_121 = _io_exe_rd_10_resp_T_120 | _io_exe_rd_10_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_122 = _io_exe_rd_10_resp_T_121 | _io_exe_rd_10_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_123 = _io_exe_rd_10_resp_T_122 | _io_exe_rd_10_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_124 = _io_exe_rd_10_resp_T_123 | _io_exe_rd_10_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_125 = _io_exe_rd_10_resp_T_124 | _io_exe_rd_10_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_126 = _io_exe_rd_10_resp_T_125 | _io_exe_rd_10_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_127 = _io_exe_rd_10_resp_T_126 | _io_exe_rd_10_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_128 = _io_exe_rd_10_resp_T_127 | _io_exe_rd_10_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_129 = _io_exe_rd_10_resp_T_128 | _io_exe_rd_10_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_130 = _io_exe_rd_10_resp_T_129 | _io_exe_rd_10_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_131 = _io_exe_rd_10_resp_T_130 | _io_exe_rd_10_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_132 = _io_exe_rd_10_resp_T_131 | _io_exe_rd_10_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_133 = _io_exe_rd_10_resp_T_132 | _io_exe_rd_10_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_134 = _io_exe_rd_10_resp_T_133 | _io_exe_rd_10_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_10_resp_T_135 = _io_exe_rd_10_resp_T_134 | _io_exe_rd_10_resp_T_85; // @[Mux.scala 27:72]
  wire [63:0] _io_exe_rd_11_resp_T = 64'h1 << io_exe_rd_11_req_idx; // @[OneHot.scala 58:35]
  wire [31:0] _io_exe_rd_11_resp_T_52 = _io_exe_rd_11_resp_T[0] ? reg_type1_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_53 = _io_exe_rd_11_resp_T[1] ? reg_type1_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_54 = _io_exe_rd_11_resp_T[2] ? reg_type1_data_nxt_2_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_55 = _io_exe_rd_11_resp_T[3] ? reg_type1_data_nxt_3_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_56 = _io_exe_rd_11_resp_T[4] ? reg_type2_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_57 = _io_exe_rd_11_resp_T[5] ? reg_type2_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_58 = _io_exe_rd_11_resp_T[6] ? reg_type2_data_nxt_2_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_59 = _io_exe_rd_11_resp_T[7] ? reg_type2_data_nxt_3_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_60 = _io_exe_rd_11_resp_T[8] ? reg_type3_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_61 = _io_exe_rd_11_resp_T[9] ? reg_type3_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_62 = _io_exe_rd_11_resp_T[10] ? reg_type4_data_nxt_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_63 = _io_exe_rd_11_resp_T[11] ? reg_type4_data_nxt_1_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_64 = _io_exe_rd_11_resp_T[12] ? reg_type4_data_nxt_2_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_65 = _io_exe_rd_11_resp_T[13] ? reg_type4_data_nxt_3_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_66 = _io_exe_rd_11_resp_T[14] ? reg_type5_data_nxt__2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_67 = _io_exe_rd_11_resp_T[15] ? reg_type5_data_nxt_1_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_68 = _io_exe_rd_11_resp_T[16] ? reg_type5_data_nxt_2_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_69 = _io_exe_rd_11_resp_T[17] ? reg_type5_data_nxt_3_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_70 = _io_exe_rd_11_resp_T[18] ? reg_type5_data_nxt_4_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_71 = _io_exe_rd_11_resp_T[19] ? reg_type5_data_nxt_5_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_72 = _io_exe_rd_11_resp_T[20] ? reg_type5_data_nxt_6_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_73 = _io_exe_rd_11_resp_T[21] ? reg_type5_data_nxt_7_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_74 = _io_exe_rd_11_resp_T[22] ? reg_type5_data_nxt_8_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_75 = _io_exe_rd_11_resp_T[23] ? reg_type5_data_nxt_9_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_76 = _io_exe_rd_11_resp_T[24] ? reg_type5_data_nxt_10_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_77 = _io_exe_rd_11_resp_T[25] ? reg_type5_data_nxt_11_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_78 = _io_exe_rd_11_resp_T[26] ? reg_type5_data_nxt_12_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_79 = _io_exe_rd_11_resp_T[27] ? reg_type5_data_nxt_13_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_80 = _io_exe_rd_11_resp_T[28] ? reg_type5_data_nxt_14_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_81 = _io_exe_rd_11_resp_T[29] ? reg_type5_data_nxt_15_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_82 = _io_exe_rd_11_resp_T[30] ? reg_type5_data_nxt_16_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_83 = _io_exe_rd_11_resp_T[31] ? reg_type5_data_nxt_17_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_84 = _io_exe_rd_11_resp_T[32] ? reg_type5_data_nxt_18_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_85 = _io_exe_rd_11_resp_T[33] ? reg_type5_data_nxt_19_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_86 = _io_exe_rd_11_resp_T[34] ? reg_type5_data_nxt_20_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_103 = _io_exe_rd_11_resp_T_52 | _io_exe_rd_11_resp_T_53; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_104 = _io_exe_rd_11_resp_T_103 | _io_exe_rd_11_resp_T_54; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_105 = _io_exe_rd_11_resp_T_104 | _io_exe_rd_11_resp_T_55; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_106 = _io_exe_rd_11_resp_T_105 | _io_exe_rd_11_resp_T_56; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_107 = _io_exe_rd_11_resp_T_106 | _io_exe_rd_11_resp_T_57; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_108 = _io_exe_rd_11_resp_T_107 | _io_exe_rd_11_resp_T_58; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_109 = _io_exe_rd_11_resp_T_108 | _io_exe_rd_11_resp_T_59; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_110 = _io_exe_rd_11_resp_T_109 | _io_exe_rd_11_resp_T_60; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_111 = _io_exe_rd_11_resp_T_110 | _io_exe_rd_11_resp_T_61; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_112 = _io_exe_rd_11_resp_T_111 | _io_exe_rd_11_resp_T_62; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_113 = _io_exe_rd_11_resp_T_112 | _io_exe_rd_11_resp_T_63; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_114 = _io_exe_rd_11_resp_T_113 | _io_exe_rd_11_resp_T_64; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_115 = _io_exe_rd_11_resp_T_114 | _io_exe_rd_11_resp_T_65; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_116 = _io_exe_rd_11_resp_T_115 | _io_exe_rd_11_resp_T_66; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_117 = _io_exe_rd_11_resp_T_116 | _io_exe_rd_11_resp_T_67; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_118 = _io_exe_rd_11_resp_T_117 | _io_exe_rd_11_resp_T_68; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_119 = _io_exe_rd_11_resp_T_118 | _io_exe_rd_11_resp_T_69; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_120 = _io_exe_rd_11_resp_T_119 | _io_exe_rd_11_resp_T_70; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_121 = _io_exe_rd_11_resp_T_120 | _io_exe_rd_11_resp_T_71; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_122 = _io_exe_rd_11_resp_T_121 | _io_exe_rd_11_resp_T_72; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_123 = _io_exe_rd_11_resp_T_122 | _io_exe_rd_11_resp_T_73; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_124 = _io_exe_rd_11_resp_T_123 | _io_exe_rd_11_resp_T_74; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_125 = _io_exe_rd_11_resp_T_124 | _io_exe_rd_11_resp_T_75; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_126 = _io_exe_rd_11_resp_T_125 | _io_exe_rd_11_resp_T_76; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_127 = _io_exe_rd_11_resp_T_126 | _io_exe_rd_11_resp_T_77; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_128 = _io_exe_rd_11_resp_T_127 | _io_exe_rd_11_resp_T_78; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_129 = _io_exe_rd_11_resp_T_128 | _io_exe_rd_11_resp_T_79; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_130 = _io_exe_rd_11_resp_T_129 | _io_exe_rd_11_resp_T_80; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_131 = _io_exe_rd_11_resp_T_130 | _io_exe_rd_11_resp_T_81; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_132 = _io_exe_rd_11_resp_T_131 | _io_exe_rd_11_resp_T_82; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_133 = _io_exe_rd_11_resp_T_132 | _io_exe_rd_11_resp_T_83; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_134 = _io_exe_rd_11_resp_T_133 | _io_exe_rd_11_resp_T_84; // @[Mux.scala 27:72]
  wire [31:0] _io_exe_rd_11_resp_T_135 = _io_exe_rd_11_resp_T_134 | _io_exe_rd_11_resp_T_85; // @[Mux.scala 27:72]
  assign io_exe_rd_0_resp = _io_exe_rd_0_resp_T_151 | _io_exe_rd_0_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_1_resp = _io_exe_rd_1_resp_T_151 | _io_exe_rd_1_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_2_resp = _io_exe_rd_2_resp_T_151 | _io_exe_rd_2_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_3_resp = _io_exe_rd_3_resp_T_151 | _io_exe_rd_3_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_4_resp = _io_exe_rd_4_resp_T_151 | _io_exe_rd_4_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_5_resp = _io_exe_rd_5_resp_T_151 | _io_exe_rd_5_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_6_resp = _io_exe_rd_6_resp_T_151 | _io_exe_rd_6_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_7_resp = _io_exe_rd_7_resp_T_151 | _io_exe_rd_7_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_8_resp = _io_exe_rd_8_resp_T_151 | _io_exe_rd_8_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_9_resp = _io_exe_rd_9_resp_T_151 | _io_exe_rd_9_resp_T_102; // @[Mux.scala 27:72]
  assign io_exe_rd_10_resp = _io_exe_rd_10_resp_T_135 | _io_exe_rd_10_resp_T_86; // @[Mux.scala 27:72]
  assign io_exe_rd_11_resp = _io_exe_rd_11_resp_T_135 | _io_exe_rd_11_resp_T_86; // @[Mux.scala 27:72]
  assign io_dec_rd_0 = reg_type2_data_2_0; // @[regfile.scala 150:16]
  assign io_dec_rd_1 = reg_type2_data_3_0; // @[regfile.scala 151:16]
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type1_data_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h0) begin
      reg_type1_data_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h0) begin
      reg_type1_data_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h0) begin
      reg_type1_data_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h0) begin
      reg_type1_data_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type1_data_0 <= _GEN_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type1_data_1_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1) begin
      reg_type1_data_1_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1) begin
      reg_type1_data_1_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1) begin
      reg_type1_data_1_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1) begin
      reg_type1_data_1_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type1_data_1_0 <= _GEN_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type1_data_2_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h2) begin
      reg_type1_data_2_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h2) begin
      reg_type1_data_2_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h2) begin
      reg_type1_data_2_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h2) begin
      reg_type1_data_2_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type1_data_2_0 <= _GEN_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type1_data_3_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h3) begin
      reg_type1_data_3_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h3) begin
      reg_type1_data_3_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h3) begin
      reg_type1_data_3_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h3) begin
      reg_type1_data_3_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type1_data_3_0 <= _GEN_19;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type2_data_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h4) begin
      reg_type2_data_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h4) begin
      reg_type2_data_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h4) begin
      reg_type2_data_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h4) begin
      reg_type2_data_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type2_data_0 <= _GEN_30;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type2_data_1_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h5) begin
      reg_type2_data_1_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h5) begin
      reg_type2_data_1_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h5) begin
      reg_type2_data_1_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h5) begin
      reg_type2_data_1_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type2_data_1_0 <= _GEN_41;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type2_data_2_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h6) begin
      reg_type2_data_2_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h6) begin
      reg_type2_data_2_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h6) begin
      reg_type2_data_2_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h6) begin
      reg_type2_data_2_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type2_data_2_0 <= _GEN_52;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type2_data_3_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h7) begin
      reg_type2_data_3_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h7) begin
      reg_type2_data_3_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h7) begin
      reg_type2_data_3_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h7) begin
      reg_type2_data_3_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type2_data_3_0 <= _GEN_63;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type3_data_0 <= 32'h800000;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h8) begin
      reg_type3_data_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h8) begin
      reg_type3_data_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h8) begin
      reg_type3_data_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h8) begin
      reg_type3_data_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type3_data_0 <= _GEN_69;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type3_data_1_0 <= 32'h800000;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h9) begin
      reg_type3_data_1_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h9) begin
      reg_type3_data_1_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h9) begin
      reg_type3_data_1_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h9) begin
      reg_type3_data_1_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type3_data_1_0 <= _GEN_75;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type4_data_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'ha) begin
      reg_type4_data_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'ha) begin
      reg_type4_data_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'ha) begin
      reg_type4_data_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'ha) begin
      reg_type4_data_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type4_data_0 <= _GEN_81;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type4_data_1_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hb) begin
      reg_type4_data_1_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hb) begin
      reg_type4_data_1_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hb) begin
      reg_type4_data_1_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hb) begin
      reg_type4_data_1_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type4_data_1_0 <= _GEN_87;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type4_data_2_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hc) begin
      reg_type4_data_2_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hc) begin
      reg_type4_data_2_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hc) begin
      reg_type4_data_2_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hc) begin
      reg_type4_data_2_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type4_data_2_0 <= _GEN_93;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type4_data_3_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hd) begin
      reg_type4_data_3_0 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hd) begin
      reg_type4_data_3_0 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hd) begin
      reg_type4_data_3_0 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hd) begin
      reg_type4_data_3_0 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type4_data_3_0 <= _GEN_99;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data__0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he) begin
      reg_type5_data__0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he) begin
      reg_type5_data__0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he) begin
      reg_type5_data__0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he) begin
      reg_type5_data__0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data__0 <= _GEN_108;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data__1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he) begin
      reg_type5_data__1 <= reg_type5_data__0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he) begin
      reg_type5_data__1 <= reg_type5_data__0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he) begin
      reg_type5_data__1 <= reg_type5_data__0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he) begin
      reg_type5_data__1 <= reg_type5_data__0;
    end else begin
      reg_type5_data__1 <= _GEN_109;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data__2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he) begin
      reg_type5_data__2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he) begin
      reg_type5_data__2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he) begin
      reg_type5_data__2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he) begin
      reg_type5_data__2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data__2 <= _GEN_110;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data__3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'he) begin
      reg_type5_data__3 <= reg_type5_data__2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'he) begin
      reg_type5_data__3 <= reg_type5_data__2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'he) begin
      reg_type5_data__3 <= reg_type5_data__2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'he) begin
      reg_type5_data__3 <= reg_type5_data__2;
    end else begin
      reg_type5_data__3 <= _GEN_111;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_1_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf) begin
      reg_type5_data_1_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf) begin
      reg_type5_data_1_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf) begin
      reg_type5_data_1_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf) begin
      reg_type5_data_1_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_1_0 <= _GEN_132;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_1_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf) begin
      reg_type5_data_1_1 <= reg_type5_data_1_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf) begin
      reg_type5_data_1_1 <= reg_type5_data_1_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf) begin
      reg_type5_data_1_1 <= reg_type5_data_1_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf) begin
      reg_type5_data_1_1 <= reg_type5_data_1_0;
    end else begin
      reg_type5_data_1_1 <= _GEN_133;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_1_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf) begin
      reg_type5_data_1_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf) begin
      reg_type5_data_1_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf) begin
      reg_type5_data_1_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf) begin
      reg_type5_data_1_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_1_2 <= _GEN_134;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_1_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'hf) begin
      reg_type5_data_1_3 <= reg_type5_data_1_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'hf) begin
      reg_type5_data_1_3 <= reg_type5_data_1_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'hf) begin
      reg_type5_data_1_3 <= reg_type5_data_1_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'hf) begin
      reg_type5_data_1_3 <= reg_type5_data_1_2;
    end else begin
      reg_type5_data_1_3 <= _GEN_135;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_2_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10) begin
      reg_type5_data_2_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10) begin
      reg_type5_data_2_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10) begin
      reg_type5_data_2_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10) begin
      reg_type5_data_2_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_2_0 <= _GEN_156;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_2_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10) begin
      reg_type5_data_2_1 <= reg_type5_data_2_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10) begin
      reg_type5_data_2_1 <= reg_type5_data_2_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10) begin
      reg_type5_data_2_1 <= reg_type5_data_2_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10) begin
      reg_type5_data_2_1 <= reg_type5_data_2_0;
    end else begin
      reg_type5_data_2_1 <= _GEN_157;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_2_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10) begin
      reg_type5_data_2_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10) begin
      reg_type5_data_2_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10) begin
      reg_type5_data_2_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10) begin
      reg_type5_data_2_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_2_2 <= _GEN_158;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_2_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h10) begin
      reg_type5_data_2_3 <= reg_type5_data_2_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h10) begin
      reg_type5_data_2_3 <= reg_type5_data_2_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h10) begin
      reg_type5_data_2_3 <= reg_type5_data_2_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h10) begin
      reg_type5_data_2_3 <= reg_type5_data_2_2;
    end else begin
      reg_type5_data_2_3 <= _GEN_159;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_3_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11) begin
      reg_type5_data_3_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11) begin
      reg_type5_data_3_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11) begin
      reg_type5_data_3_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11) begin
      reg_type5_data_3_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_3_0 <= _GEN_180;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_3_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11) begin
      reg_type5_data_3_1 <= reg_type5_data_3_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11) begin
      reg_type5_data_3_1 <= reg_type5_data_3_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11) begin
      reg_type5_data_3_1 <= reg_type5_data_3_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11) begin
      reg_type5_data_3_1 <= reg_type5_data_3_0;
    end else begin
      reg_type5_data_3_1 <= _GEN_181;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_3_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11) begin
      reg_type5_data_3_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11) begin
      reg_type5_data_3_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11) begin
      reg_type5_data_3_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11) begin
      reg_type5_data_3_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_3_2 <= _GEN_182;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_3_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h11) begin
      reg_type5_data_3_3 <= reg_type5_data_3_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h11) begin
      reg_type5_data_3_3 <= reg_type5_data_3_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h11) begin
      reg_type5_data_3_3 <= reg_type5_data_3_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h11) begin
      reg_type5_data_3_3 <= reg_type5_data_3_2;
    end else begin
      reg_type5_data_3_3 <= _GEN_183;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_4_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12) begin
      reg_type5_data_4_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12) begin
      reg_type5_data_4_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12) begin
      reg_type5_data_4_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12) begin
      reg_type5_data_4_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_4_0 <= _GEN_204;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_4_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12) begin
      reg_type5_data_4_1 <= reg_type5_data_4_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12) begin
      reg_type5_data_4_1 <= reg_type5_data_4_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12) begin
      reg_type5_data_4_1 <= reg_type5_data_4_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12) begin
      reg_type5_data_4_1 <= reg_type5_data_4_0;
    end else begin
      reg_type5_data_4_1 <= _GEN_205;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_4_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12) begin
      reg_type5_data_4_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12) begin
      reg_type5_data_4_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12) begin
      reg_type5_data_4_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12) begin
      reg_type5_data_4_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_4_2 <= _GEN_206;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_4_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h12) begin
      reg_type5_data_4_3 <= reg_type5_data_4_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h12) begin
      reg_type5_data_4_3 <= reg_type5_data_4_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h12) begin
      reg_type5_data_4_3 <= reg_type5_data_4_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h12) begin
      reg_type5_data_4_3 <= reg_type5_data_4_2;
    end else begin
      reg_type5_data_4_3 <= _GEN_207;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_5_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13) begin
      reg_type5_data_5_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13) begin
      reg_type5_data_5_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13) begin
      reg_type5_data_5_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13) begin
      reg_type5_data_5_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_5_0 <= _GEN_228;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_5_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13) begin
      reg_type5_data_5_1 <= reg_type5_data_5_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13) begin
      reg_type5_data_5_1 <= reg_type5_data_5_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13) begin
      reg_type5_data_5_1 <= reg_type5_data_5_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13) begin
      reg_type5_data_5_1 <= reg_type5_data_5_0;
    end else begin
      reg_type5_data_5_1 <= _GEN_229;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_5_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13) begin
      reg_type5_data_5_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13) begin
      reg_type5_data_5_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13) begin
      reg_type5_data_5_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13) begin
      reg_type5_data_5_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_5_2 <= _GEN_230;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_5_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h13) begin
      reg_type5_data_5_3 <= reg_type5_data_5_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h13) begin
      reg_type5_data_5_3 <= reg_type5_data_5_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h13) begin
      reg_type5_data_5_3 <= reg_type5_data_5_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h13) begin
      reg_type5_data_5_3 <= reg_type5_data_5_2;
    end else begin
      reg_type5_data_5_3 <= _GEN_231;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_6_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14) begin
      reg_type5_data_6_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14) begin
      reg_type5_data_6_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14) begin
      reg_type5_data_6_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14) begin
      reg_type5_data_6_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_6_0 <= _GEN_252;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_6_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14) begin
      reg_type5_data_6_1 <= reg_type5_data_6_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14) begin
      reg_type5_data_6_1 <= reg_type5_data_6_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14) begin
      reg_type5_data_6_1 <= reg_type5_data_6_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14) begin
      reg_type5_data_6_1 <= reg_type5_data_6_0;
    end else begin
      reg_type5_data_6_1 <= _GEN_253;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_6_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14) begin
      reg_type5_data_6_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14) begin
      reg_type5_data_6_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14) begin
      reg_type5_data_6_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14) begin
      reg_type5_data_6_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_6_2 <= _GEN_254;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_6_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h14) begin
      reg_type5_data_6_3 <= reg_type5_data_6_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h14) begin
      reg_type5_data_6_3 <= reg_type5_data_6_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h14) begin
      reg_type5_data_6_3 <= reg_type5_data_6_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h14) begin
      reg_type5_data_6_3 <= reg_type5_data_6_2;
    end else begin
      reg_type5_data_6_3 <= _GEN_255;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_7_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15) begin
      reg_type5_data_7_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15) begin
      reg_type5_data_7_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15) begin
      reg_type5_data_7_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15) begin
      reg_type5_data_7_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_7_0 <= _GEN_276;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_7_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15) begin
      reg_type5_data_7_1 <= reg_type5_data_7_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15) begin
      reg_type5_data_7_1 <= reg_type5_data_7_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15) begin
      reg_type5_data_7_1 <= reg_type5_data_7_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15) begin
      reg_type5_data_7_1 <= reg_type5_data_7_0;
    end else begin
      reg_type5_data_7_1 <= _GEN_277;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_7_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15) begin
      reg_type5_data_7_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15) begin
      reg_type5_data_7_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15) begin
      reg_type5_data_7_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15) begin
      reg_type5_data_7_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_7_2 <= _GEN_278;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_7_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h15) begin
      reg_type5_data_7_3 <= reg_type5_data_7_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h15) begin
      reg_type5_data_7_3 <= reg_type5_data_7_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h15) begin
      reg_type5_data_7_3 <= reg_type5_data_7_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h15) begin
      reg_type5_data_7_3 <= reg_type5_data_7_2;
    end else begin
      reg_type5_data_7_3 <= _GEN_279;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_8_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16) begin
      reg_type5_data_8_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16) begin
      reg_type5_data_8_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16) begin
      reg_type5_data_8_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16) begin
      reg_type5_data_8_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_8_0 <= _GEN_300;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_8_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16) begin
      reg_type5_data_8_1 <= reg_type5_data_8_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16) begin
      reg_type5_data_8_1 <= reg_type5_data_8_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16) begin
      reg_type5_data_8_1 <= reg_type5_data_8_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16) begin
      reg_type5_data_8_1 <= reg_type5_data_8_0;
    end else begin
      reg_type5_data_8_1 <= _GEN_301;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_8_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16) begin
      reg_type5_data_8_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16) begin
      reg_type5_data_8_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16) begin
      reg_type5_data_8_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16) begin
      reg_type5_data_8_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_8_2 <= _GEN_302;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_8_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h16) begin
      reg_type5_data_8_3 <= reg_type5_data_8_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h16) begin
      reg_type5_data_8_3 <= reg_type5_data_8_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h16) begin
      reg_type5_data_8_3 <= reg_type5_data_8_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h16) begin
      reg_type5_data_8_3 <= reg_type5_data_8_2;
    end else begin
      reg_type5_data_8_3 <= _GEN_303;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_9_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17) begin
      reg_type5_data_9_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17) begin
      reg_type5_data_9_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17) begin
      reg_type5_data_9_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17) begin
      reg_type5_data_9_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_9_0 <= _GEN_324;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_9_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17) begin
      reg_type5_data_9_1 <= reg_type5_data_9_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17) begin
      reg_type5_data_9_1 <= reg_type5_data_9_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17) begin
      reg_type5_data_9_1 <= reg_type5_data_9_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17) begin
      reg_type5_data_9_1 <= reg_type5_data_9_0;
    end else begin
      reg_type5_data_9_1 <= _GEN_325;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_9_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17) begin
      reg_type5_data_9_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17) begin
      reg_type5_data_9_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17) begin
      reg_type5_data_9_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17) begin
      reg_type5_data_9_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_9_2 <= _GEN_326;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_9_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h17) begin
      reg_type5_data_9_3 <= reg_type5_data_9_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h17) begin
      reg_type5_data_9_3 <= reg_type5_data_9_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h17) begin
      reg_type5_data_9_3 <= reg_type5_data_9_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h17) begin
      reg_type5_data_9_3 <= reg_type5_data_9_2;
    end else begin
      reg_type5_data_9_3 <= _GEN_327;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_10_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18) begin
      reg_type5_data_10_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18) begin
      reg_type5_data_10_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18) begin
      reg_type5_data_10_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18) begin
      reg_type5_data_10_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_10_0 <= _GEN_348;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_10_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18) begin
      reg_type5_data_10_1 <= reg_type5_data_10_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18) begin
      reg_type5_data_10_1 <= reg_type5_data_10_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18) begin
      reg_type5_data_10_1 <= reg_type5_data_10_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18) begin
      reg_type5_data_10_1 <= reg_type5_data_10_0;
    end else begin
      reg_type5_data_10_1 <= _GEN_349;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_10_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18) begin
      reg_type5_data_10_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18) begin
      reg_type5_data_10_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18) begin
      reg_type5_data_10_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18) begin
      reg_type5_data_10_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_10_2 <= _GEN_350;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_10_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h18) begin
      reg_type5_data_10_3 <= reg_type5_data_10_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h18) begin
      reg_type5_data_10_3 <= reg_type5_data_10_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h18) begin
      reg_type5_data_10_3 <= reg_type5_data_10_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h18) begin
      reg_type5_data_10_3 <= reg_type5_data_10_2;
    end else begin
      reg_type5_data_10_3 <= _GEN_351;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_11_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19) begin
      reg_type5_data_11_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19) begin
      reg_type5_data_11_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19) begin
      reg_type5_data_11_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19) begin
      reg_type5_data_11_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_11_0 <= _GEN_372;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_11_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19) begin
      reg_type5_data_11_1 <= reg_type5_data_11_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19) begin
      reg_type5_data_11_1 <= reg_type5_data_11_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19) begin
      reg_type5_data_11_1 <= reg_type5_data_11_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19) begin
      reg_type5_data_11_1 <= reg_type5_data_11_0;
    end else begin
      reg_type5_data_11_1 <= _GEN_373;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_11_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19) begin
      reg_type5_data_11_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19) begin
      reg_type5_data_11_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19) begin
      reg_type5_data_11_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19) begin
      reg_type5_data_11_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_11_2 <= _GEN_374;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_11_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h19) begin
      reg_type5_data_11_3 <= reg_type5_data_11_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h19) begin
      reg_type5_data_11_3 <= reg_type5_data_11_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h19) begin
      reg_type5_data_11_3 <= reg_type5_data_11_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h19) begin
      reg_type5_data_11_3 <= reg_type5_data_11_2;
    end else begin
      reg_type5_data_11_3 <= _GEN_375;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_12_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a) begin
      reg_type5_data_12_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a) begin
      reg_type5_data_12_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a) begin
      reg_type5_data_12_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a) begin
      reg_type5_data_12_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_12_0 <= _GEN_396;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_12_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a) begin
      reg_type5_data_12_1 <= reg_type5_data_12_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a) begin
      reg_type5_data_12_1 <= reg_type5_data_12_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a) begin
      reg_type5_data_12_1 <= reg_type5_data_12_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a) begin
      reg_type5_data_12_1 <= reg_type5_data_12_0;
    end else begin
      reg_type5_data_12_1 <= _GEN_397;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_12_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a) begin
      reg_type5_data_12_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a) begin
      reg_type5_data_12_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a) begin
      reg_type5_data_12_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a) begin
      reg_type5_data_12_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_12_2 <= _GEN_398;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_12_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1a) begin
      reg_type5_data_12_3 <= reg_type5_data_12_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1a) begin
      reg_type5_data_12_3 <= reg_type5_data_12_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1a) begin
      reg_type5_data_12_3 <= reg_type5_data_12_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1a) begin
      reg_type5_data_12_3 <= reg_type5_data_12_2;
    end else begin
      reg_type5_data_12_3 <= _GEN_399;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_13_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b) begin
      reg_type5_data_13_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b) begin
      reg_type5_data_13_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b) begin
      reg_type5_data_13_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b) begin
      reg_type5_data_13_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_13_0 <= _GEN_420;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_13_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b) begin
      reg_type5_data_13_1 <= reg_type5_data_13_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b) begin
      reg_type5_data_13_1 <= reg_type5_data_13_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b) begin
      reg_type5_data_13_1 <= reg_type5_data_13_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b) begin
      reg_type5_data_13_1 <= reg_type5_data_13_0;
    end else begin
      reg_type5_data_13_1 <= _GEN_421;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_13_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b) begin
      reg_type5_data_13_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b) begin
      reg_type5_data_13_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b) begin
      reg_type5_data_13_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b) begin
      reg_type5_data_13_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_13_2 <= _GEN_422;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_13_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1b) begin
      reg_type5_data_13_3 <= reg_type5_data_13_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1b) begin
      reg_type5_data_13_3 <= reg_type5_data_13_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1b) begin
      reg_type5_data_13_3 <= reg_type5_data_13_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1b) begin
      reg_type5_data_13_3 <= reg_type5_data_13_2;
    end else begin
      reg_type5_data_13_3 <= _GEN_423;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_14_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c) begin
      reg_type5_data_14_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c) begin
      reg_type5_data_14_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c) begin
      reg_type5_data_14_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c) begin
      reg_type5_data_14_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_14_0 <= _GEN_444;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_14_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c) begin
      reg_type5_data_14_1 <= reg_type5_data_14_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c) begin
      reg_type5_data_14_1 <= reg_type5_data_14_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c) begin
      reg_type5_data_14_1 <= reg_type5_data_14_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c) begin
      reg_type5_data_14_1 <= reg_type5_data_14_0;
    end else begin
      reg_type5_data_14_1 <= _GEN_445;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_14_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c) begin
      reg_type5_data_14_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c) begin
      reg_type5_data_14_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c) begin
      reg_type5_data_14_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c) begin
      reg_type5_data_14_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_14_2 <= _GEN_446;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_14_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1c) begin
      reg_type5_data_14_3 <= reg_type5_data_14_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1c) begin
      reg_type5_data_14_3 <= reg_type5_data_14_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1c) begin
      reg_type5_data_14_3 <= reg_type5_data_14_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1c) begin
      reg_type5_data_14_3 <= reg_type5_data_14_2;
    end else begin
      reg_type5_data_14_3 <= _GEN_447;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_15_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d) begin
      reg_type5_data_15_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d) begin
      reg_type5_data_15_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d) begin
      reg_type5_data_15_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d) begin
      reg_type5_data_15_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_15_0 <= _GEN_468;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_15_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d) begin
      reg_type5_data_15_1 <= reg_type5_data_15_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d) begin
      reg_type5_data_15_1 <= reg_type5_data_15_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d) begin
      reg_type5_data_15_1 <= reg_type5_data_15_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d) begin
      reg_type5_data_15_1 <= reg_type5_data_15_0;
    end else begin
      reg_type5_data_15_1 <= _GEN_469;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_15_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d) begin
      reg_type5_data_15_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d) begin
      reg_type5_data_15_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d) begin
      reg_type5_data_15_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d) begin
      reg_type5_data_15_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_15_2 <= _GEN_470;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_15_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1d) begin
      reg_type5_data_15_3 <= reg_type5_data_15_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1d) begin
      reg_type5_data_15_3 <= reg_type5_data_15_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1d) begin
      reg_type5_data_15_3 <= reg_type5_data_15_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1d) begin
      reg_type5_data_15_3 <= reg_type5_data_15_2;
    end else begin
      reg_type5_data_15_3 <= _GEN_471;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_16_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e) begin
      reg_type5_data_16_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e) begin
      reg_type5_data_16_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e) begin
      reg_type5_data_16_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e) begin
      reg_type5_data_16_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_16_0 <= _GEN_492;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_16_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e) begin
      reg_type5_data_16_1 <= reg_type5_data_16_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e) begin
      reg_type5_data_16_1 <= reg_type5_data_16_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e) begin
      reg_type5_data_16_1 <= reg_type5_data_16_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e) begin
      reg_type5_data_16_1 <= reg_type5_data_16_0;
    end else begin
      reg_type5_data_16_1 <= _GEN_493;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_16_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e) begin
      reg_type5_data_16_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e) begin
      reg_type5_data_16_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e) begin
      reg_type5_data_16_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e) begin
      reg_type5_data_16_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_16_2 <= _GEN_494;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_16_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1e) begin
      reg_type5_data_16_3 <= reg_type5_data_16_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1e) begin
      reg_type5_data_16_3 <= reg_type5_data_16_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1e) begin
      reg_type5_data_16_3 <= reg_type5_data_16_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1e) begin
      reg_type5_data_16_3 <= reg_type5_data_16_2;
    end else begin
      reg_type5_data_16_3 <= _GEN_495;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_17_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f) begin
      reg_type5_data_17_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f) begin
      reg_type5_data_17_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f) begin
      reg_type5_data_17_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f) begin
      reg_type5_data_17_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_17_0 <= _GEN_516;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_17_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f) begin
      reg_type5_data_17_1 <= reg_type5_data_17_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f) begin
      reg_type5_data_17_1 <= reg_type5_data_17_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f) begin
      reg_type5_data_17_1 <= reg_type5_data_17_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f) begin
      reg_type5_data_17_1 <= reg_type5_data_17_0;
    end else begin
      reg_type5_data_17_1 <= _GEN_517;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_17_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f) begin
      reg_type5_data_17_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f) begin
      reg_type5_data_17_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f) begin
      reg_type5_data_17_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f) begin
      reg_type5_data_17_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_17_2 <= _GEN_518;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_17_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h1f) begin
      reg_type5_data_17_3 <= reg_type5_data_17_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h1f) begin
      reg_type5_data_17_3 <= reg_type5_data_17_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h1f) begin
      reg_type5_data_17_3 <= reg_type5_data_17_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h1f) begin
      reg_type5_data_17_3 <= reg_type5_data_17_2;
    end else begin
      reg_type5_data_17_3 <= _GEN_519;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_18_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20) begin
      reg_type5_data_18_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20) begin
      reg_type5_data_18_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20) begin
      reg_type5_data_18_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20) begin
      reg_type5_data_18_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_18_0 <= _GEN_540;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_18_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20) begin
      reg_type5_data_18_1 <= reg_type5_data_18_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20) begin
      reg_type5_data_18_1 <= reg_type5_data_18_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20) begin
      reg_type5_data_18_1 <= reg_type5_data_18_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20) begin
      reg_type5_data_18_1 <= reg_type5_data_18_0;
    end else begin
      reg_type5_data_18_1 <= _GEN_541;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_18_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20) begin
      reg_type5_data_18_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20) begin
      reg_type5_data_18_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20) begin
      reg_type5_data_18_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20) begin
      reg_type5_data_18_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_18_2 <= _GEN_542;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_18_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h20) begin
      reg_type5_data_18_3 <= reg_type5_data_18_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h20) begin
      reg_type5_data_18_3 <= reg_type5_data_18_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h20) begin
      reg_type5_data_18_3 <= reg_type5_data_18_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h20) begin
      reg_type5_data_18_3 <= reg_type5_data_18_2;
    end else begin
      reg_type5_data_18_3 <= _GEN_543;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_19_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21) begin
      reg_type5_data_19_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21) begin
      reg_type5_data_19_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21) begin
      reg_type5_data_19_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21) begin
      reg_type5_data_19_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_19_0 <= _GEN_564;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_19_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21) begin
      reg_type5_data_19_1 <= reg_type5_data_19_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21) begin
      reg_type5_data_19_1 <= reg_type5_data_19_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21) begin
      reg_type5_data_19_1 <= reg_type5_data_19_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21) begin
      reg_type5_data_19_1 <= reg_type5_data_19_0;
    end else begin
      reg_type5_data_19_1 <= _GEN_565;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_19_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21) begin
      reg_type5_data_19_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21) begin
      reg_type5_data_19_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21) begin
      reg_type5_data_19_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21) begin
      reg_type5_data_19_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_19_2 <= _GEN_566;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_19_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h21) begin
      reg_type5_data_19_3 <= reg_type5_data_19_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h21) begin
      reg_type5_data_19_3 <= reg_type5_data_19_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h21) begin
      reg_type5_data_19_3 <= reg_type5_data_19_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h21) begin
      reg_type5_data_19_3 <= reg_type5_data_19_2;
    end else begin
      reg_type5_data_19_3 <= _GEN_567;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_20_0 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22) begin
      reg_type5_data_20_0 <= 32'h0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22) begin
      reg_type5_data_20_0 <= io_exe_wb_4_wdata1;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22) begin
      reg_type5_data_20_0 <= io_exe_wb_3_wdata1;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22) begin
      reg_type5_data_20_0 <= io_exe_wb_2_wdata1;
    end else begin
      reg_type5_data_20_0 <= _GEN_588;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_20_1 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22) begin
      reg_type5_data_20_1 <= reg_type5_data_20_0;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22) begin
      reg_type5_data_20_1 <= reg_type5_data_20_0;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22) begin
      reg_type5_data_20_1 <= reg_type5_data_20_0;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22) begin
      reg_type5_data_20_1 <= reg_type5_data_20_0;
    end else begin
      reg_type5_data_20_1 <= _GEN_589;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_20_2 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22) begin
      reg_type5_data_20_2 <= io_exe_wb_5_wdata2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22) begin
      reg_type5_data_20_2 <= io_exe_wb_4_wdata2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22) begin
      reg_type5_data_20_2 <= io_exe_wb_3_wdata2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22) begin
      reg_type5_data_20_2 <= io_exe_wb_2_wdata2;
    end else begin
      reg_type5_data_20_2 <= _GEN_590;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      reg_type5_data_20_3 <= 32'h0;
    end else if (io_exe_wb_5_vld & io_exe_wb_5_gregidx == 6'h22) begin
      reg_type5_data_20_3 <= reg_type5_data_20_2;
    end else if (io_exe_wb_4_vld & io_exe_wb_4_gregidx == 6'h22) begin
      reg_type5_data_20_3 <= reg_type5_data_20_2;
    end else if (io_exe_wb_3_vld & io_exe_wb_3_gregidx == 6'h22) begin
      reg_type5_data_20_3 <= reg_type5_data_20_2;
    end else if (io_exe_wb_2_vld & io_exe_wb_2_gregidx == 6'h22) begin
      reg_type5_data_20_3 <= reg_type5_data_20_2;
    end else begin
      reg_type5_data_20_3 <= _GEN_591;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_type1_data_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_type1_data_1_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_type1_data_2_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_type1_data_3_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_type2_data_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_type2_data_1_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_type2_data_2_0 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_type2_data_3_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_type3_data_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_type3_data_1_0 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_type4_data_0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_type4_data_1_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_type4_data_2_0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_type4_data_3_0 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_type5_data__0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_type5_data__1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_type5_data__2 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_type5_data__3 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_type5_data_1_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_type5_data_1_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_type5_data_1_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_type5_data_1_3 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_type5_data_2_0 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_type5_data_2_1 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_type5_data_2_2 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_type5_data_2_3 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_type5_data_3_0 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_type5_data_3_1 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_type5_data_3_2 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_type5_data_3_3 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_type5_data_4_0 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_type5_data_4_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  reg_type5_data_4_2 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  reg_type5_data_4_3 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  reg_type5_data_5_0 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  reg_type5_data_5_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  reg_type5_data_5_2 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_type5_data_5_3 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  reg_type5_data_6_0 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  reg_type5_data_6_1 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  reg_type5_data_6_2 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  reg_type5_data_6_3 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  reg_type5_data_7_0 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  reg_type5_data_7_1 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  reg_type5_data_7_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  reg_type5_data_7_3 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  reg_type5_data_8_0 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  reg_type5_data_8_1 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  reg_type5_data_8_2 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  reg_type5_data_8_3 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  reg_type5_data_9_0 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  reg_type5_data_9_1 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  reg_type5_data_9_2 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  reg_type5_data_9_3 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  reg_type5_data_10_0 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  reg_type5_data_10_1 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  reg_type5_data_10_2 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  reg_type5_data_10_3 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  reg_type5_data_11_0 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  reg_type5_data_11_1 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  reg_type5_data_11_2 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  reg_type5_data_11_3 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  reg_type5_data_12_0 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  reg_type5_data_12_1 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  reg_type5_data_12_2 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  reg_type5_data_12_3 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  reg_type5_data_13_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  reg_type5_data_13_1 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  reg_type5_data_13_2 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  reg_type5_data_13_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  reg_type5_data_14_0 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  reg_type5_data_14_1 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  reg_type5_data_14_2 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  reg_type5_data_14_3 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  reg_type5_data_15_0 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  reg_type5_data_15_1 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  reg_type5_data_15_2 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  reg_type5_data_15_3 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  reg_type5_data_16_0 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  reg_type5_data_16_1 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  reg_type5_data_16_2 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  reg_type5_data_16_3 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  reg_type5_data_17_0 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  reg_type5_data_17_1 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  reg_type5_data_17_2 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  reg_type5_data_17_3 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  reg_type5_data_18_0 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  reg_type5_data_18_1 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  reg_type5_data_18_2 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  reg_type5_data_18_3 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  reg_type5_data_19_0 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  reg_type5_data_19_1 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  reg_type5_data_19_2 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  reg_type5_data_19_3 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  reg_type5_data_20_0 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  reg_type5_data_20_1 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  reg_type5_data_20_2 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  reg_type5_data_20_3 = _RAND_97[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    reg_type1_data_0 = 32'h0;
  end
  if (reset) begin
    reg_type1_data_1_0 = 32'h0;
  end
  if (reset) begin
    reg_type1_data_2_0 = 32'h0;
  end
  if (reset) begin
    reg_type1_data_3_0 = 32'h0;
  end
  if (reset) begin
    reg_type2_data_0 = 32'h0;
  end
  if (reset) begin
    reg_type2_data_1_0 = 32'h0;
  end
  if (reset) begin
    reg_type2_data_2_0 = 32'h0;
  end
  if (reset) begin
    reg_type2_data_3_0 = 32'h0;
  end
  if (reset) begin
    reg_type3_data_0 = 32'h800000;
  end
  if (reset) begin
    reg_type3_data_1_0 = 32'h800000;
  end
  if (reset) begin
    reg_type4_data_0 = 32'h0;
  end
  if (reset) begin
    reg_type4_data_1_0 = 32'h0;
  end
  if (reset) begin
    reg_type4_data_2_0 = 32'h0;
  end
  if (reset) begin
    reg_type4_data_3_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data__0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data__1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data__2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data__3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_1_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_1_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_1_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_1_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_2_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_2_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_2_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_2_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_3_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_3_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_3_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_3_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_4_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_4_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_4_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_4_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_5_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_5_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_5_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_5_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_6_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_6_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_6_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_6_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_7_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_7_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_7_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_7_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_8_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_8_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_8_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_8_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_9_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_9_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_9_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_9_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_10_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_10_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_10_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_10_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_11_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_11_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_11_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_11_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_12_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_12_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_12_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_12_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_13_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_13_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_13_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_13_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_14_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_14_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_14_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_14_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_15_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_15_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_15_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_15_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_16_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_16_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_16_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_16_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_17_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_17_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_17_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_17_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_18_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_18_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_18_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_18_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_19_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_19_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_19_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_19_3 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_20_0 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_20_1 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_20_2 = 32'h0;
  end
  if (reset) begin
    reg_type5_data_20_3 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MacUnit(
  input         clock,
  input         reset,
  output        io_uopin_ready,
  input         io_uopin_valid,
  input  [2:0]  io_uopin_bits_vlen,
  input         io_uopin_bits_select,
  input         io_uopin_bits_drc,
  input         io_uopin_bits_pow,
  input         io_uopin_bits_loop,
  input         io_uopin_bits_drcgain,
  input         io_uopin_bits_drcnum,
  input         io_uopin_bits_srcreq_0_valid,
  input         io_uopin_bits_srcreq_0_isgroup,
  input         io_uopin_bits_srcreq_0_iscoef,
  input  [5:0]  io_uopin_bits_srcreq_0_idx,
  input         io_uopin_bits_srcreq_0_busy,
  input         io_uopin_bits_srcreq_0_wkupidx_0,
  input         io_uopin_bits_srcreq_0_wkupidx_1,
  input         io_uopin_bits_srcreq_0_wkupidx_2,
  input         io_uopin_bits_srcreq_0_wkupidx_3,
  input         io_uopin_bits_srcreq_0_wkupidx_4,
  input         io_uopin_bits_srcreq_0_wkupidx_5,
  input         io_uopin_bits_srcreq_1_valid,
  input         io_uopin_bits_srcreq_1_isgroup,
  input         io_uopin_bits_srcreq_1_iscoef,
  input  [5:0]  io_uopin_bits_srcreq_1_idx,
  input         io_uopin_bits_srcreq_1_busy,
  input         io_uopin_bits_srcreq_1_wkupidx_0,
  input         io_uopin_bits_srcreq_1_wkupidx_1,
  input         io_uopin_bits_srcreq_1_wkupidx_2,
  input         io_uopin_bits_srcreq_1_wkupidx_3,
  input         io_uopin_bits_srcreq_1_wkupidx_4,
  input         io_uopin_bits_srcreq_1_wkupidx_5,
  input         io_uopin_bits_srcreq_2_valid,
  input         io_uopin_bits_srcreq_2_isgroup,
  input         io_uopin_bits_srcreq_2_iscoef,
  input  [5:0]  io_uopin_bits_srcreq_2_idx,
  input         io_uopin_bits_srcreq_2_busy,
  input         io_uopin_bits_srcreq_2_wkupidx_0,
  input         io_uopin_bits_srcreq_2_wkupidx_1,
  input         io_uopin_bits_srcreq_2_wkupidx_2,
  input         io_uopin_bits_srcreq_2_wkupidx_3,
  input         io_uopin_bits_srcreq_2_wkupidx_4,
  input         io_uopin_bits_srcreq_2_wkupidx_5,
  input         io_uopin_bits_srcreq_3_valid,
  input         io_uopin_bits_srcreq_3_isgroup,
  input         io_uopin_bits_srcreq_3_iscoef,
  input  [5:0]  io_uopin_bits_srcreq_3_idx,
  input         io_uopin_bits_srcreq_3_busy,
  input         io_uopin_bits_srcreq_3_wkupidx_0,
  input         io_uopin_bits_srcreq_3_wkupidx_1,
  input         io_uopin_bits_srcreq_3_wkupidx_2,
  input         io_uopin_bits_srcreq_3_wkupidx_3,
  input         io_uopin_bits_srcreq_3_wkupidx_4,
  input         io_uopin_bits_srcreq_3_wkupidx_5,
  input         io_uopin_bits_srcreq_4_valid,
  input         io_uopin_bits_srcreq_4_isgroup,
  input         io_uopin_bits_srcreq_4_iscoef,
  input  [5:0]  io_uopin_bits_srcreq_4_idx,
  input         io_uopin_bits_srcreq_4_busy,
  input         io_uopin_bits_srcreq_4_wkupidx_0,
  input         io_uopin_bits_srcreq_4_wkupidx_1,
  input         io_uopin_bits_srcreq_4_wkupidx_2,
  input         io_uopin_bits_srcreq_4_wkupidx_3,
  input         io_uopin_bits_srcreq_4_wkupidx_4,
  input         io_uopin_bits_srcreq_4_wkupidx_5,
  input         io_uopin_bits_srcreq_5_valid,
  input         io_uopin_bits_srcreq_5_isgroup,
  input         io_uopin_bits_srcreq_5_iscoef,
  input  [5:0]  io_uopin_bits_srcreq_5_idx,
  input         io_uopin_bits_srcreq_5_busy,
  input         io_uopin_bits_srcreq_5_wkupidx_0,
  input         io_uopin_bits_srcreq_5_wkupidx_1,
  input         io_uopin_bits_srcreq_5_wkupidx_2,
  input         io_uopin_bits_srcreq_5_wkupidx_3,
  input         io_uopin_bits_srcreq_5_wkupidx_4,
  input         io_uopin_bits_srcreq_5_wkupidx_5,
  input         io_uopin_bits_wbvld,
  input  [5:0]  io_uopin_bits_wbreq,
  input         io_uopin_bits_waridx_0,
  input         io_uopin_bits_waridx_1,
  input         io_uopin_bits_waridx_2,
  input         io_uopin_bits_waridx_3,
  input         io_uopin_bits_waridx_4,
  input         io_uopin_bits_wawidx_0,
  input         io_uopin_bits_wawidx_1,
  input         io_uopin_bits_wawidx_2,
  input         io_uopin_bits_wawidx_3,
  input         io_uopin_bits_wawidx_4,
  output        io_rfreq_0_req_isgroup,
  output        io_rfreq_0_req_iscoef,
  output [5:0]  io_rfreq_0_req_idx,
  output [2:0]  io_rfreq_0_req_gidx,
  input  [31:0] io_rfreq_0_resp,
  output        io_rfreq_1_req_isgroup,
  output        io_rfreq_1_req_iscoef,
  output [5:0]  io_rfreq_1_req_idx,
  output [2:0]  io_rfreq_1_req_gidx,
  output        io_rfreq_1_req_sel,
  input  [31:0] io_rfreq_1_resp,
  output [31:0] io_wbreq_wdata1,
  output [31:0] io_wbreq_wdata2,
  output        io_wbreq_vld,
  output [5:0]  io_wbreq_gregidx,
  output        io_fwd_wkup_valid,
  output [5:0]  io_fwd_wkup_bits,
  output        io_empty,
  input         io_raw_wkup_0_valid,
  input  [5:0]  io_raw_wkup_0_bits,
  input         io_raw_wkup_1_valid,
  input  [5:0]  io_raw_wkup_1_bits,
  input         io_raw_wkup_2_valid,
  input  [5:0]  io_raw_wkup_2_bits,
  input         io_raw_wkup_3_valid,
  input  [5:0]  io_raw_wkup_3_bits,
  input         io_raw_wkup_4_valid,
  input  [5:0]  io_raw_wkup_4_bits,
  input         io_raw_wkup_5_valid,
  input  [5:0]  io_raw_wkup_5_bits,
  output        io_wbcheck_valid,
  output [5:0]  io_wbcheck_bits,
  output        io_r_check_0_valid,
  output [5:0]  io_r_check_0_bits,
  output        io_r_check_1_valid,
  output [5:0]  io_r_check_1_bits,
  output        io_r_check_2_valid,
  output [5:0]  io_r_check_2_bits,
  output        io_r_check_3_valid,
  output [5:0]  io_r_check_3_bits,
  output        io_r_check_4_valid,
  output [5:0]  io_r_check_4_bits,
  output        io_r_check_5_valid,
  output [5:0]  io_r_check_5_bits,
  input         io_other_flop_0,
  input         io_other_flop_1,
  input         io_other_flop_2,
  input         io_other_flop_3,
  input         io_other_flop_4,
  output        io_flop,
  input  [31:0] io_coef_subch_drc_th,
  input  [31:0] io_coef_subch_drc_offset,
  input         io_coef_subch_drc_drcen,
  input         io_coef_mainch_ch0_autoloop,
  input  [31:0] io_coef_mainch_drc_th,
  input  [31:0] io_coef_mainch_drc_offset,
  input         io_coef_mainch_drc_drcen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
`endif // RANDOMIZE_REG_INIT
  reg  s1_uop_valid; // @[macu.scala 26:23]
  reg [2:0] s1_uop_bits_vlen; // @[macu.scala 26:23]
  reg  s1_uop_bits_select; // @[macu.scala 26:23]
  reg  s1_uop_bits_drc; // @[macu.scala 26:23]
  reg  s1_uop_bits_pow; // @[macu.scala 26:23]
  reg  s1_uop_bits_loop; // @[macu.scala 26:23]
  reg  s1_uop_bits_drcgain; // @[macu.scala 26:23]
  reg  s1_uop_bits_drcnum; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_valid; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_isgroup; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_iscoef; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_srcreq_0_idx; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_busy; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_wkupidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_wkupidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_wkupidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_wkupidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_wkupidx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_0_wkupidx_5; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_valid; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_isgroup; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_iscoef; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_srcreq_1_idx; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_busy; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_wkupidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_wkupidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_wkupidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_wkupidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_wkupidx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_1_wkupidx_5; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_valid; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_isgroup; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_iscoef; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_srcreq_2_idx; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_busy; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_wkupidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_wkupidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_wkupidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_wkupidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_wkupidx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_2_wkupidx_5; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_valid; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_isgroup; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_iscoef; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_srcreq_3_idx; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_busy; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_wkupidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_wkupidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_wkupidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_wkupidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_wkupidx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_3_wkupidx_5; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_valid; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_isgroup; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_iscoef; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_srcreq_4_idx; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_busy; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_wkupidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_wkupidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_wkupidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_wkupidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_wkupidx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_4_wkupidx_5; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_valid; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_isgroup; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_iscoef; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_srcreq_5_idx; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_busy; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_wkupidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_wkupidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_wkupidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_wkupidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_wkupidx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_srcreq_5_wkupidx_5; // @[macu.scala 26:23]
  reg  s1_uop_bits_wbvld; // @[macu.scala 26:23]
  reg [5:0] s1_uop_bits_wbreq; // @[macu.scala 26:23]
  reg  s1_uop_bits_waridx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_waridx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_waridx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_waridx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_waridx_4; // @[macu.scala 26:23]
  reg  s1_uop_bits_wawidx_0; // @[macu.scala 26:23]
  reg  s1_uop_bits_wawidx_1; // @[macu.scala 26:23]
  reg  s1_uop_bits_wawidx_2; // @[macu.scala 26:23]
  reg  s1_uop_bits_wawidx_3; // @[macu.scala 26:23]
  reg  s1_uop_bits_wawidx_4; // @[macu.scala 26:23]
  reg [1:0] s1_state; // @[macu.scala 30:25]
  reg  s2_vld; // @[macu.scala 33:24]
  reg  s2_wb; // @[macu.scala 34:24]
  reg [5:0] s2_wbidx; // @[macu.scala 35:24]
  reg [31:0] s2_data_0; // @[macu.scala 38:24]
  reg [31:0] s2_data_1; // @[macu.scala 38:24]
  reg [31:0] s2_data_2; // @[macu.scala 38:24]
  wire  _no_depd_T_7 = s1_uop_bits_wawidx_0 | s1_uop_bits_wawidx_1 | s1_uop_bits_wawidx_2 | s1_uop_bits_wawidx_3 |
    s1_uop_bits_wawidx_4; // @[macu.scala 43:47]
  wire  no_depd = ~(s1_uop_bits_waridx_0 | s1_uop_bits_waridx_1 | s1_uop_bits_waridx_2 | s1_uop_bits_waridx_3 |
    s1_uop_bits_waridx_4 | _no_depd_T_7); // @[macu.scala 42:17]
  wire  _T = s1_state == 2'h2; // @[macu.scala 80:18]
  wire  _GEN_204 = 3'h1 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_1_valid : s1_uop_bits_srcreq_0_valid; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_205 = 3'h2 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_2_valid : _GEN_204; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_206 = 3'h3 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_3_valid : _GEN_205; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_207 = 3'h4 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_4_valid : _GEN_206; // @[macu.scala 100:13 macu.scala 100:13]
  wire  rf_req_0_valid = 3'h5 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_5_valid : _GEN_207; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_180 = 3'h1 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_1_busy : s1_uop_bits_srcreq_0_busy; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_181 = 3'h2 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_2_busy : _GEN_180; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_182 = 3'h3 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_3_busy : _GEN_181; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_183 = 3'h4 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_4_busy : _GEN_182; // @[macu.scala 100:13 macu.scala 100:13]
  wire  rf_req_0_busy = 3'h5 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_5_busy : _GEN_183; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _req2_idx_T = s1_state == 2'h1; // @[macu.scala 95:31]
  wire [2:0] _req2_idx_T_2 = s1_uop_bits_vlen + 3'h1; // @[macu.scala 95:57]
  wire [2:0] req2_idx = s1_state == 2'h1 ? _req2_idx_T_2 : 3'h5; // @[macu.scala 95:21]
  wire  _GEN_138 = 3'h1 == req2_idx ? s1_uop_bits_srcreq_1_valid : s1_uop_bits_srcreq_0_valid; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_139 = 3'h2 == req2_idx ? s1_uop_bits_srcreq_2_valid : _GEN_138; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_140 = 3'h3 == req2_idx ? s1_uop_bits_srcreq_3_valid : _GEN_139; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_141 = 3'h4 == req2_idx ? s1_uop_bits_srcreq_4_valid : _GEN_140; // @[macu.scala 99:13 macu.scala 99:13]
  wire  rf_req_1_valid = 3'h5 == req2_idx ? s1_uop_bits_srcreq_5_valid : _GEN_141; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_114 = 3'h1 == req2_idx ? s1_uop_bits_srcreq_1_busy : s1_uop_bits_srcreq_0_busy; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_115 = 3'h2 == req2_idx ? s1_uop_bits_srcreq_2_busy : _GEN_114; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_116 = 3'h3 == req2_idx ? s1_uop_bits_srcreq_3_busy : _GEN_115; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_117 = 3'h4 == req2_idx ? s1_uop_bits_srcreq_4_busy : _GEN_116; // @[macu.scala 99:13 macu.scala 99:13]
  wire  rf_req_1_busy = 3'h5 == req2_idx ? s1_uop_bits_srcreq_5_busy : _GEN_117; // @[macu.scala 99:13 macu.scala 99:13]
  wire  read_en = (rf_req_0_valid & ~rf_req_0_busy | ~rf_req_0_valid) & (rf_req_1_valid & ~rf_req_1_busy | ~
    rf_req_1_valid) & s1_uop_valid; // @[macu.scala 114:75]
  wire  _T_1 = s1_state == 2'h2 & read_en; // @[macu.scala 80:28]
  wire [2:0] _s1_uop_bits_vlen_T_1 = s1_uop_bits_vlen - 3'h1; // @[macu.scala 81:42]
  wire  _T_5 = s1_state == 2'h3; // @[macu.scala 85:60]
  wire  out__0 = s1_uop_bits_wawidx_0 & ~io_other_flop_0; // @[macu.scala 64:41]
  wire  out__1 = s1_uop_bits_wawidx_1 & ~io_other_flop_1; // @[macu.scala 64:41]
  wire  out__2 = s1_uop_bits_wawidx_2 & ~io_other_flop_2; // @[macu.scala 64:41]
  wire  out__3 = s1_uop_bits_wawidx_3 & ~io_other_flop_3; // @[macu.scala 64:41]
  wire  out__4 = s1_uop_bits_wawidx_4 & ~io_other_flop_4; // @[macu.scala 64:41]
  wire  out_1_0 = s1_uop_bits_waridx_0 & ~io_other_flop_0; // @[macu.scala 64:41]
  wire  out_1_1 = s1_uop_bits_waridx_1 & ~io_other_flop_1; // @[macu.scala 64:41]
  wire  out_1_2 = s1_uop_bits_waridx_2 & ~io_other_flop_2; // @[macu.scala 64:41]
  wire  out_1_3 = s1_uop_bits_waridx_3 & ~io_other_flop_3; // @[macu.scala 64:41]
  wire  out_1_4 = s1_uop_bits_waridx_4 & ~io_other_flop_4; // @[macu.scala 64:41]
  wire [7:0] _T_27 = 8'h1 << s1_uop_bits_vlen; // @[OneHot.scala 58:35]
  wire [7:0] _T_28 = 8'h1 << req2_idx; // @[OneHot.scala 58:35]
  wire [7:0] _T_29 = _T_27 | _T_28; // @[macu.scala 101:43]
  wire  read_vec_0 = _T_29[0]; // @[macu.scala 101:77]
  wire  _s1_uop_bits_srcreq_0_out_valid_T_1 = ~(read_vec_0 & read_en); // @[macu.scala 51:33]
  wire  s1_uop_bits_srcreq_0_out_valid = s1_uop_bits_srcreq_0_valid & ~(read_vec_0 & read_en); // @[macu.scala 51:30]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_0_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_0_out_wkupidx_0_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_0 = s1_uop_bits_srcreq_0_wkupidx_0 & _s1_uop_bits_srcreq_0_out_wkupidx_0_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_0_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_0_out_wkupidx_1_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_1 = s1_uop_bits_srcreq_0_wkupidx_1 & _s1_uop_bits_srcreq_0_out_wkupidx_1_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_0_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_0_out_wkupidx_2_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_2 = s1_uop_bits_srcreq_0_wkupidx_2 & _s1_uop_bits_srcreq_0_out_wkupidx_2_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_0_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_0_out_wkupidx_3_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_3 = s1_uop_bits_srcreq_0_wkupidx_3 & _s1_uop_bits_srcreq_0_out_wkupidx_3_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_0_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_0_out_wkupidx_4_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_4 = s1_uop_bits_srcreq_0_wkupidx_4 & _s1_uop_bits_srcreq_0_out_wkupidx_4_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_0_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_0_out_wkupidx_5_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_5 = s1_uop_bits_srcreq_0_wkupidx_5 & _s1_uop_bits_srcreq_0_out_wkupidx_5_T_2; // @[macu.scala 54:40]
  wire  s1_uop_bits_srcreq_0_out_busy = s1_uop_bits_srcreq_0_out_wkupidx_0 | s1_uop_bits_srcreq_0_out_wkupidx_1 |
    s1_uop_bits_srcreq_0_out_wkupidx_2 | s1_uop_bits_srcreq_0_out_wkupidx_3 | s1_uop_bits_srcreq_0_out_wkupidx_4 |
    s1_uop_bits_srcreq_0_out_wkupidx_5; // @[macu.scala 58:37]
  wire  read_vec_1 = _T_29[1]; // @[macu.scala 101:77]
  wire  _s1_uop_bits_srcreq_1_out_valid_T_1 = ~(read_vec_1 & read_en); // @[macu.scala 51:33]
  wire  s1_uop_bits_srcreq_1_out_valid = s1_uop_bits_srcreq_1_valid & ~(read_vec_1 & read_en); // @[macu.scala 51:30]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_1_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_1_out_wkupidx_0_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_0 = s1_uop_bits_srcreq_1_wkupidx_0 & _s1_uop_bits_srcreq_1_out_wkupidx_0_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_1_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_1_out_wkupidx_1_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_1 = s1_uop_bits_srcreq_1_wkupidx_1 & _s1_uop_bits_srcreq_1_out_wkupidx_1_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_1_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_1_out_wkupidx_2_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_2 = s1_uop_bits_srcreq_1_wkupidx_2 & _s1_uop_bits_srcreq_1_out_wkupidx_2_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_1_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_1_out_wkupidx_3_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_3 = s1_uop_bits_srcreq_1_wkupidx_3 & _s1_uop_bits_srcreq_1_out_wkupidx_3_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_1_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_1_out_wkupidx_4_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_4 = s1_uop_bits_srcreq_1_wkupidx_4 & _s1_uop_bits_srcreq_1_out_wkupidx_4_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_1_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_1_out_wkupidx_5_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_5 = s1_uop_bits_srcreq_1_wkupidx_5 & _s1_uop_bits_srcreq_1_out_wkupidx_5_T_2; // @[macu.scala 54:40]
  wire  s1_uop_bits_srcreq_1_out_busy = s1_uop_bits_srcreq_1_out_wkupidx_0 | s1_uop_bits_srcreq_1_out_wkupidx_1 |
    s1_uop_bits_srcreq_1_out_wkupidx_2 | s1_uop_bits_srcreq_1_out_wkupidx_3 | s1_uop_bits_srcreq_1_out_wkupidx_4 |
    s1_uop_bits_srcreq_1_out_wkupidx_5; // @[macu.scala 58:37]
  wire  read_vec_2 = _T_29[2]; // @[macu.scala 101:77]
  wire  _s1_uop_bits_srcreq_2_out_valid_T_1 = ~(read_vec_2 & read_en); // @[macu.scala 51:33]
  wire  s1_uop_bits_srcreq_2_out_valid = s1_uop_bits_srcreq_2_valid & ~(read_vec_2 & read_en); // @[macu.scala 51:30]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_2_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_2_out_wkupidx_0_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_2_out_wkupidx_0 = s1_uop_bits_srcreq_2_wkupidx_0 & _s1_uop_bits_srcreq_2_out_wkupidx_0_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_2_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_2_out_wkupidx_1_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_2_out_wkupidx_1 = s1_uop_bits_srcreq_2_wkupidx_1 & _s1_uop_bits_srcreq_2_out_wkupidx_1_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_2_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_2_out_wkupidx_2_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_2_out_wkupidx_2 = s1_uop_bits_srcreq_2_wkupidx_2 & _s1_uop_bits_srcreq_2_out_wkupidx_2_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_2_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_2_out_wkupidx_3_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_2_out_wkupidx_3 = s1_uop_bits_srcreq_2_wkupidx_3 & _s1_uop_bits_srcreq_2_out_wkupidx_3_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_2_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_2_out_wkupidx_4_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_2_out_wkupidx_4 = s1_uop_bits_srcreq_2_wkupidx_4 & _s1_uop_bits_srcreq_2_out_wkupidx_4_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_2_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_2_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_2_out_wkupidx_5_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_2_out_wkupidx_5 = s1_uop_bits_srcreq_2_wkupidx_5 & _s1_uop_bits_srcreq_2_out_wkupidx_5_T_2; // @[macu.scala 54:40]
  wire  s1_uop_bits_srcreq_2_out_busy = s1_uop_bits_srcreq_2_out_wkupidx_0 | s1_uop_bits_srcreq_2_out_wkupidx_1 |
    s1_uop_bits_srcreq_2_out_wkupidx_2 | s1_uop_bits_srcreq_2_out_wkupidx_3 | s1_uop_bits_srcreq_2_out_wkupidx_4 |
    s1_uop_bits_srcreq_2_out_wkupidx_5; // @[macu.scala 58:37]
  wire  read_vec_3 = _T_29[3]; // @[macu.scala 101:77]
  wire  _s1_uop_bits_srcreq_3_out_valid_T_1 = ~(read_vec_3 & read_en); // @[macu.scala 51:33]
  wire  s1_uop_bits_srcreq_3_out_valid = s1_uop_bits_srcreq_3_valid & ~(read_vec_3 & read_en); // @[macu.scala 51:30]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_3_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_3_out_wkupidx_0_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_3_out_wkupidx_0 = s1_uop_bits_srcreq_3_wkupidx_0 & _s1_uop_bits_srcreq_3_out_wkupidx_0_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_3_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_3_out_wkupidx_1_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_3_out_wkupidx_1 = s1_uop_bits_srcreq_3_wkupidx_1 & _s1_uop_bits_srcreq_3_out_wkupidx_1_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_3_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_3_out_wkupidx_2_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_3_out_wkupidx_2 = s1_uop_bits_srcreq_3_wkupidx_2 & _s1_uop_bits_srcreq_3_out_wkupidx_2_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_3_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_3_out_wkupidx_3_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_3_out_wkupidx_3 = s1_uop_bits_srcreq_3_wkupidx_3 & _s1_uop_bits_srcreq_3_out_wkupidx_3_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_3_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_3_out_wkupidx_4_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_3_out_wkupidx_4 = s1_uop_bits_srcreq_3_wkupidx_4 & _s1_uop_bits_srcreq_3_out_wkupidx_4_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_3_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_3_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_3_out_wkupidx_5_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_3_out_wkupidx_5 = s1_uop_bits_srcreq_3_wkupidx_5 & _s1_uop_bits_srcreq_3_out_wkupidx_5_T_2; // @[macu.scala 54:40]
  wire  s1_uop_bits_srcreq_3_out_busy = s1_uop_bits_srcreq_3_out_wkupidx_0 | s1_uop_bits_srcreq_3_out_wkupidx_1 |
    s1_uop_bits_srcreq_3_out_wkupidx_2 | s1_uop_bits_srcreq_3_out_wkupidx_3 | s1_uop_bits_srcreq_3_out_wkupidx_4 |
    s1_uop_bits_srcreq_3_out_wkupidx_5; // @[macu.scala 58:37]
  wire  read_vec_4 = _T_29[4]; // @[macu.scala 101:77]
  wire  _s1_uop_bits_srcreq_4_out_valid_T_1 = ~(read_vec_4 & read_en); // @[macu.scala 51:33]
  wire  s1_uop_bits_srcreq_4_out_valid = s1_uop_bits_srcreq_4_valid & ~(read_vec_4 & read_en); // @[macu.scala 51:30]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_4_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_4_out_wkupidx_0_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_4_out_wkupidx_0 = s1_uop_bits_srcreq_4_wkupidx_0 & _s1_uop_bits_srcreq_4_out_wkupidx_0_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_4_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_4_out_wkupidx_1_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_4_out_wkupidx_1 = s1_uop_bits_srcreq_4_wkupidx_1 & _s1_uop_bits_srcreq_4_out_wkupidx_1_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_4_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_4_out_wkupidx_2_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_4_out_wkupidx_2 = s1_uop_bits_srcreq_4_wkupidx_2 & _s1_uop_bits_srcreq_4_out_wkupidx_2_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_4_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_4_out_wkupidx_3_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_4_out_wkupidx_3 = s1_uop_bits_srcreq_4_wkupidx_3 & _s1_uop_bits_srcreq_4_out_wkupidx_3_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_4_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_4_out_wkupidx_4_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_4_out_wkupidx_4 = s1_uop_bits_srcreq_4_wkupidx_4 & _s1_uop_bits_srcreq_4_out_wkupidx_4_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_4_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_4_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_4_out_wkupidx_5_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_4_out_wkupidx_5 = s1_uop_bits_srcreq_4_wkupidx_5 & _s1_uop_bits_srcreq_4_out_wkupidx_5_T_2; // @[macu.scala 54:40]
  wire  s1_uop_bits_srcreq_4_out_busy = s1_uop_bits_srcreq_4_out_wkupidx_0 | s1_uop_bits_srcreq_4_out_wkupidx_1 |
    s1_uop_bits_srcreq_4_out_wkupidx_2 | s1_uop_bits_srcreq_4_out_wkupidx_3 | s1_uop_bits_srcreq_4_out_wkupidx_4 |
    s1_uop_bits_srcreq_4_out_wkupidx_5; // @[macu.scala 58:37]
  wire  read_vec_5 = _T_29[5]; // @[macu.scala 101:77]
  wire  _s1_uop_bits_srcreq_5_out_valid_T = read_vec_5 & read_en; // @[macu.scala 49:41]
  wire  _s1_uop_bits_srcreq_5_out_valid_T_1 = s1_uop_bits_vlen == 3'h0; // @[macu.scala 49:73]
  wire  s1_uop_bits_srcreq_5_out_valid = s1_uop_bits_srcreq_5_valid & ~(read_vec_5 & read_en & s1_uop_bits_vlen == 3'h0)
    ; // @[macu.scala 49:30]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_5_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_5_out_wkupidx_0_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_5_out_wkupidx_0 = s1_uop_bits_srcreq_5_wkupidx_0 & _s1_uop_bits_srcreq_5_out_wkupidx_0_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_5_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_5_out_wkupidx_1_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_5_out_wkupidx_1 = s1_uop_bits_srcreq_5_wkupidx_1 & _s1_uop_bits_srcreq_5_out_wkupidx_1_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_5_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_5_out_wkupidx_2_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_5_out_wkupidx_2 = s1_uop_bits_srcreq_5_wkupidx_2 & _s1_uop_bits_srcreq_5_out_wkupidx_2_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_5_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_5_out_wkupidx_3_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_5_out_wkupidx_3 = s1_uop_bits_srcreq_5_wkupidx_3 & _s1_uop_bits_srcreq_5_out_wkupidx_3_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_5_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_5_out_wkupidx_4_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_5_out_wkupidx_4 = s1_uop_bits_srcreq_5_wkupidx_4 & _s1_uop_bits_srcreq_5_out_wkupidx_4_T_2; // @[macu.scala 54:40]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_5_idx; // @[macu.scala 56:51]
  wire  _s1_uop_bits_srcreq_5_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_5_out_wkupidx_5_T_1; // @[macu.scala 55:52]
  wire  s1_uop_bits_srcreq_5_out_wkupidx_5 = s1_uop_bits_srcreq_5_wkupidx_5 & _s1_uop_bits_srcreq_5_out_wkupidx_5_T_2; // @[macu.scala 54:40]
  wire  s1_uop_bits_srcreq_5_out_busy = s1_uop_bits_srcreq_5_out_wkupidx_0 | s1_uop_bits_srcreq_5_out_wkupidx_1 |
    s1_uop_bits_srcreq_5_out_wkupidx_2 | s1_uop_bits_srcreq_5_out_wkupidx_3 | s1_uop_bits_srcreq_5_out_wkupidx_4 |
    s1_uop_bits_srcreq_5_out_wkupidx_5; // @[macu.scala 58:37]
  reg  select; // @[macu.scala 96:23]
  wire [31:0] data_diff = io_rfreq_0_resp - io_rfreq_1_resp; // @[macu.scala 97:36]
  wire [5:0] _GEN_120 = 3'h1 == req2_idx ? s1_uop_bits_srcreq_1_idx : s1_uop_bits_srcreq_0_idx; // @[macu.scala 99:13 macu.scala 99:13]
  wire [5:0] _GEN_121 = 3'h2 == req2_idx ? s1_uop_bits_srcreq_2_idx : _GEN_120; // @[macu.scala 99:13 macu.scala 99:13]
  wire [5:0] _GEN_122 = 3'h3 == req2_idx ? s1_uop_bits_srcreq_3_idx : _GEN_121; // @[macu.scala 99:13 macu.scala 99:13]
  wire [5:0] _GEN_123 = 3'h4 == req2_idx ? s1_uop_bits_srcreq_4_idx : _GEN_122; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_126 = 3'h1 == req2_idx ? s1_uop_bits_srcreq_1_iscoef : s1_uop_bits_srcreq_0_iscoef; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_127 = 3'h2 == req2_idx ? s1_uop_bits_srcreq_2_iscoef : _GEN_126; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_128 = 3'h3 == req2_idx ? s1_uop_bits_srcreq_3_iscoef : _GEN_127; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_129 = 3'h4 == req2_idx ? s1_uop_bits_srcreq_4_iscoef : _GEN_128; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_132 = 3'h1 == req2_idx ? s1_uop_bits_srcreq_1_isgroup : s1_uop_bits_srcreq_0_isgroup; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_133 = 3'h2 == req2_idx ? s1_uop_bits_srcreq_2_isgroup : _GEN_132; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_134 = 3'h3 == req2_idx ? s1_uop_bits_srcreq_3_isgroup : _GEN_133; // @[macu.scala 99:13 macu.scala 99:13]
  wire  _GEN_135 = 3'h4 == req2_idx ? s1_uop_bits_srcreq_4_isgroup : _GEN_134; // @[macu.scala 99:13 macu.scala 99:13]
  wire [5:0] _GEN_186 = 3'h1 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_1_idx : s1_uop_bits_srcreq_0_idx; // @[macu.scala 100:13 macu.scala 100:13]
  wire [5:0] _GEN_187 = 3'h2 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_2_idx : _GEN_186; // @[macu.scala 100:13 macu.scala 100:13]
  wire [5:0] _GEN_188 = 3'h3 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_3_idx : _GEN_187; // @[macu.scala 100:13 macu.scala 100:13]
  wire [5:0] _GEN_189 = 3'h4 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_4_idx : _GEN_188; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_192 = 3'h1 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_1_iscoef : s1_uop_bits_srcreq_0_iscoef; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_193 = 3'h2 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_2_iscoef : _GEN_192; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_194 = 3'h3 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_3_iscoef : _GEN_193; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_195 = 3'h4 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_4_iscoef : _GEN_194; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_198 = 3'h1 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_1_isgroup : s1_uop_bits_srcreq_0_isgroup; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_199 = 3'h2 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_2_isgroup : _GEN_198; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_200 = 3'h3 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_3_isgroup : _GEN_199; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _GEN_201 = 3'h4 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_4_isgroup : _GEN_200; // @[macu.scala 100:13 macu.scala 100:13]
  wire  _select_T_1 = _req2_idx_T & read_en; // @[macu.scala 102:35]
  wire [1:0] idle_nxt = io_uopin_bits_select | io_uopin_bits_loop ? 2'h1 : 2'h2; // @[macu.scala 115:21]
  wire  _T_37 = s1_state == 2'h0; // @[macu.scala 120:17]
  wire  _s1_nxt_state_T = io_uopin_ready & io_uopin_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _s1_nxt_state_T_1 = _s1_nxt_state_T ? idle_nxt : 2'h0; // @[macu.scala 121:24]
  wire [1:0] _s1_nxt_state_T_2 = read_en ? 2'h2 : 2'h1; // @[macu.scala 124:24]
  wire [1:0] _s1_nxt_state_T_5 = no_depd ? _s1_nxt_state_T_1 : 2'h3; // @[macu.scala 127:26]
  wire [1:0] _GEN_209 = _s1_uop_bits_srcreq_5_out_valid_T_1 & read_en ? _s1_nxt_state_T_5 : s1_state; // @[macu.scala 126:49 macu.scala 127:20 macu.scala 119:16]
  wire [1:0] _GEN_210 = _T_5 ? _s1_nxt_state_T_5 : s1_state; // @[macu.scala 131:34 macu.scala 132:18 macu.scala 119:16]
  wire [1:0] _GEN_211 = _T ? _GEN_209 : _GEN_210; // @[macu.scala 125:33]
  wire [1:0] _GEN_212 = _req2_idx_T ? _s1_nxt_state_T_2 : _GEN_211; // @[macu.scala 123:33 macu.scala 124:18]
  wire [1:0] s1_nxt_state = s1_state == 2'h0 ? _s1_nxt_state_T_1 : _GEN_212; // @[macu.scala 120:28 macu.scala 121:18]
  wire  _io_flop_T_1 = _T_5 & no_depd; // @[macu.scala 137:35]
  wire  _io_flop_T_7 = _T_1 & read_en & _s1_uop_bits_srcreq_5_out_valid_T_1 & no_depd; // @[macu.scala 138:77]
  wire  flop = _T_1 & no_depd & _s1_uop_bits_srcreq_5_out_valid_T_1 | _io_flop_T_1; // @[macu.scala 140:86]
  reg [31:0] loop_data; // @[macu.scala 157:26]
  wire  drc1 = ~s1_uop_bits_drcnum; // @[macu.scala 158:17]
  wire [31:0] drccoef_th = drc1 ? io_coef_mainch_drc_th : io_coef_subch_drc_th; // @[macu.scala 159:20]
  wire  drccoef_drcen = drc1 ? io_coef_mainch_drc_drcen : io_coef_subch_drc_drcen; // @[macu.scala 159:20]
  wire [31:0] _drc_data_T_1 = io_rfreq_0_resp - drccoef_th; // @[macu.scala 160:41]
  reg  start; // @[macu.scala 166:22]
  wire  _GEN_214 = start & read_en & _T ? 1'h0 : start; // @[macu.scala 170:54 macu.scala 171:11 macu.scala 166:22]
  wire [31:0] _s1_data_0_out_T_1 = 32'sh0 - $signed(io_rfreq_0_resp); // @[macu.scala 72:46]
  wire [31:0] s1_data_0_out = io_rfreq_0_resp[31] ? _s1_data_0_out_T_1 : io_rfreq_0_resp; // @[macu.scala 72:15]
  wire [63:0] _product_T_2 = $signed(s2_data_0) * $signed(s2_data_1); // @[macu.scala 206:54]
  wire [40:0] _GEN_301 = _product_T_2[63:23];
  wire [31:0] product = _GEN_301[31:0];
  wire [31:0] _s2_dout_T_1 = s2_vld ? $signed(product) : $signed(32'sh0); // @[macu.scala 207:18]
  wire [31:0] s2_dout = $signed(_s2_dout_T_1) + $signed(s2_data_2); // @[macu.scala 207:71]
  reg  io_fwd_wkup_valid_REG; // @[macu.scala 198:40]
  reg  io_wbreq_vld_REG; // @[macu.scala 212:26]
  reg [5:0] io_wbreq_gregidx_REG; // @[macu.scala 213:30]
  reg [31:0] io_wbreq_wdata1_REG; // @[macu.scala 214:29]
  reg [31:0] io_wbreq_wdata2_REG; // @[macu.scala 215:29]
  assign io_uopin_ready = flop | _T_37; // @[macu.scala 154:26]
  assign io_rfreq_0_req_isgroup = 3'h5 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_5_isgroup : _GEN_201; // @[macu.scala 100:13 macu.scala 100:13]
  assign io_rfreq_0_req_iscoef = 3'h5 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_5_iscoef : _GEN_195; // @[macu.scala 100:13 macu.scala 100:13]
  assign io_rfreq_0_req_idx = 3'h5 == s1_uop_bits_vlen ? s1_uop_bits_srcreq_5_idx : _GEN_189; // @[macu.scala 100:13 macu.scala 100:13]
  assign io_rfreq_0_req_gidx = s1_uop_bits_vlen; // @[macu.scala 109:26]
  assign io_rfreq_1_req_isgroup = 3'h5 == req2_idx ? s1_uop_bits_srcreq_5_isgroup : _GEN_135; // @[macu.scala 99:13 macu.scala 99:13]
  assign io_rfreq_1_req_iscoef = 3'h5 == req2_idx ? s1_uop_bits_srcreq_5_iscoef : _GEN_129; // @[macu.scala 99:13 macu.scala 99:13]
  assign io_rfreq_1_req_idx = 3'h5 == req2_idx ? s1_uop_bits_srcreq_5_idx : _GEN_123; // @[macu.scala 99:13 macu.scala 99:13]
  assign io_rfreq_1_req_gidx = s1_uop_bits_vlen; // @[macu.scala 109:26]
  assign io_rfreq_1_req_sel = select; // @[macu.scala 112:23]
  assign io_wbreq_wdata1 = io_wbreq_wdata1_REG; // @[macu.scala 214:19]
  assign io_wbreq_wdata2 = io_wbreq_wdata2_REG; // @[macu.scala 215:19]
  assign io_wbreq_vld = io_wbreq_vld_REG; // @[macu.scala 212:16]
  assign io_wbreq_gregidx = io_wbreq_gregidx_REG; // @[macu.scala 213:20]
  assign io_fwd_wkup_valid = s2_wb & io_fwd_wkup_valid_REG; // @[macu.scala 198:30]
  assign io_fwd_wkup_bits = s2_wbidx; // @[macu.scala 199:21]
  assign io_empty = ~s1_uop_valid & ~s2_vld & ~io_wbreq_vld; // @[macu.scala 153:40]
  assign io_wbcheck_valid = s1_uop_bits_wbvld & s1_uop_valid & ~flop; // @[macu.scala 144:57]
  assign io_wbcheck_bits = s1_uop_bits_wbreq; // @[macu.scala 145:19]
  assign io_r_check_0_valid = s1_uop_valid & s1_uop_bits_srcreq_0_valid & _s1_uop_bits_srcreq_0_out_valid_T_1 & ~
    s1_uop_bits_srcreq_0_iscoef; // @[macu.scala 149:83]
  assign io_r_check_0_bits = s1_uop_bits_srcreq_0_idx; // @[macu.scala 150:25]
  assign io_r_check_1_valid = s1_uop_valid & s1_uop_bits_srcreq_1_valid & _s1_uop_bits_srcreq_1_out_valid_T_1 & ~
    s1_uop_bits_srcreq_1_iscoef; // @[macu.scala 149:83]
  assign io_r_check_1_bits = s1_uop_bits_srcreq_1_idx; // @[macu.scala 150:25]
  assign io_r_check_2_valid = s1_uop_valid & s1_uop_bits_srcreq_2_valid & _s1_uop_bits_srcreq_2_out_valid_T_1 & ~
    s1_uop_bits_srcreq_2_iscoef; // @[macu.scala 149:83]
  assign io_r_check_2_bits = s1_uop_bits_srcreq_2_idx; // @[macu.scala 150:25]
  assign io_r_check_3_valid = s1_uop_valid & s1_uop_bits_srcreq_3_valid & _s1_uop_bits_srcreq_3_out_valid_T_1 & ~
    s1_uop_bits_srcreq_3_iscoef; // @[macu.scala 149:83]
  assign io_r_check_3_bits = s1_uop_bits_srcreq_3_idx; // @[macu.scala 150:25]
  assign io_r_check_4_valid = s1_uop_valid & s1_uop_bits_srcreq_4_valid & _s1_uop_bits_srcreq_4_out_valid_T_1 & ~
    s1_uop_bits_srcreq_4_iscoef; // @[macu.scala 149:83]
  assign io_r_check_4_bits = s1_uop_bits_srcreq_4_idx; // @[macu.scala 150:25]
  assign io_r_check_5_valid = s1_uop_valid & s1_uop_bits_srcreq_5_valid & ~_s1_uop_bits_srcreq_5_out_valid_T & ~
    s1_uop_bits_srcreq_5_iscoef; // @[macu.scala 149:83]
  assign io_r_check_5_bits = s1_uop_bits_srcreq_5_idx; // @[macu.scala 150:25]
  assign io_flop = _T_5 & no_depd | _io_flop_T_7; // @[macu.scala 137:46]
  always @(posedge clock) begin
    io_fwd_wkup_valid_REG <= s1_uop_valid & s1_uop_bits_wbvld; // @[macu.scala 198:54]
    io_wbreq_vld_REG <= s2_wb; // @[macu.scala 212:26]
    io_wbreq_gregidx_REG <= s2_wbidx; // @[macu.scala 213:30]
    io_wbreq_wdata1_REG <= s2_data_0; // @[macu.scala 214:29]
    io_wbreq_wdata2_REG <= $signed(_s2_dout_T_1) + $signed(s2_data_2); // @[macu.scala 207:71]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_valid <= 1'h0;
    end else begin
      s1_uop_valid <= s1_nxt_state != 2'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_vlen <= 3'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_vlen <= io_uopin_bits_vlen;
    end else if (s1_state == 2'h2 & read_en) begin
      s1_uop_bits_vlen <= _s1_uop_bits_vlen_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_select <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_select <= io_uopin_bits_select;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_drc <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_drc <= io_uopin_bits_drc;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_pow <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_pow <= io_uopin_bits_pow;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_loop <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_loop <= io_uopin_bits_loop;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_drcgain <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_drcgain <= io_uopin_bits_drcgain;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_drcnum <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_drcnum <= io_uopin_bits_drcnum;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_valid <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_valid <= io_uopin_bits_srcreq_0_valid;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_valid <= s1_uop_bits_srcreq_0_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_isgroup <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_isgroup <= io_uopin_bits_srcreq_0_isgroup;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_iscoef <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_iscoef <= io_uopin_bits_srcreq_0_iscoef;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_idx <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_idx <= io_uopin_bits_srcreq_0_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_busy <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_busy <= io_uopin_bits_srcreq_0_busy;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_busy <= s1_uop_bits_srcreq_0_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_wkupidx_0 <= io_uopin_bits_srcreq_0_wkupidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_wkupidx_0 <= s1_uop_bits_srcreq_0_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_wkupidx_1 <= io_uopin_bits_srcreq_0_wkupidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_wkupidx_1 <= s1_uop_bits_srcreq_0_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_wkupidx_2 <= io_uopin_bits_srcreq_0_wkupidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_wkupidx_2 <= s1_uop_bits_srcreq_0_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_wkupidx_3 <= io_uopin_bits_srcreq_0_wkupidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_wkupidx_3 <= s1_uop_bits_srcreq_0_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_wkupidx_4 <= io_uopin_bits_srcreq_0_wkupidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_wkupidx_4 <= s1_uop_bits_srcreq_0_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_5 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_0_wkupidx_5 <= io_uopin_bits_srcreq_0_wkupidx_5;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_0_wkupidx_5 <= s1_uop_bits_srcreq_0_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_valid <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_valid <= io_uopin_bits_srcreq_1_valid;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_valid <= s1_uop_bits_srcreq_1_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_isgroup <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_isgroup <= io_uopin_bits_srcreq_1_isgroup;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_iscoef <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_iscoef <= io_uopin_bits_srcreq_1_iscoef;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_idx <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_idx <= io_uopin_bits_srcreq_1_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_busy <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_busy <= io_uopin_bits_srcreq_1_busy;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_busy <= s1_uop_bits_srcreq_1_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_wkupidx_0 <= io_uopin_bits_srcreq_1_wkupidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_wkupidx_0 <= s1_uop_bits_srcreq_1_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_wkupidx_1 <= io_uopin_bits_srcreq_1_wkupidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_wkupidx_1 <= s1_uop_bits_srcreq_1_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_wkupidx_2 <= io_uopin_bits_srcreq_1_wkupidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_wkupidx_2 <= s1_uop_bits_srcreq_1_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_wkupidx_3 <= io_uopin_bits_srcreq_1_wkupidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_wkupidx_3 <= s1_uop_bits_srcreq_1_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_wkupidx_4 <= io_uopin_bits_srcreq_1_wkupidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_wkupidx_4 <= s1_uop_bits_srcreq_1_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_5 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_1_wkupidx_5 <= io_uopin_bits_srcreq_1_wkupidx_5;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_1_wkupidx_5 <= s1_uop_bits_srcreq_1_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_valid <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_valid <= io_uopin_bits_srcreq_2_valid;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_valid <= s1_uop_bits_srcreq_2_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_isgroup <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_isgroup <= io_uopin_bits_srcreq_2_isgroup;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_iscoef <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_iscoef <= io_uopin_bits_srcreq_2_iscoef;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_idx <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_idx <= io_uopin_bits_srcreq_2_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_busy <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_busy <= io_uopin_bits_srcreq_2_busy;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_busy <= s1_uop_bits_srcreq_2_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_wkupidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_wkupidx_0 <= io_uopin_bits_srcreq_2_wkupidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_wkupidx_0 <= s1_uop_bits_srcreq_2_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_wkupidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_wkupidx_1 <= io_uopin_bits_srcreq_2_wkupidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_wkupidx_1 <= s1_uop_bits_srcreq_2_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_wkupidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_wkupidx_2 <= io_uopin_bits_srcreq_2_wkupidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_wkupidx_2 <= s1_uop_bits_srcreq_2_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_wkupidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_wkupidx_3 <= io_uopin_bits_srcreq_2_wkupidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_wkupidx_3 <= s1_uop_bits_srcreq_2_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_wkupidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_wkupidx_4 <= io_uopin_bits_srcreq_2_wkupidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_wkupidx_4 <= s1_uop_bits_srcreq_2_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_2_wkupidx_5 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_2_wkupidx_5 <= io_uopin_bits_srcreq_2_wkupidx_5;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_2_wkupidx_5 <= s1_uop_bits_srcreq_2_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_valid <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_valid <= io_uopin_bits_srcreq_3_valid;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_valid <= s1_uop_bits_srcreq_3_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_isgroup <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_isgroup <= io_uopin_bits_srcreq_3_isgroup;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_iscoef <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_iscoef <= io_uopin_bits_srcreq_3_iscoef;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_idx <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_idx <= io_uopin_bits_srcreq_3_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_busy <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_busy <= io_uopin_bits_srcreq_3_busy;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_busy <= s1_uop_bits_srcreq_3_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_wkupidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_wkupidx_0 <= io_uopin_bits_srcreq_3_wkupidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_wkupidx_0 <= s1_uop_bits_srcreq_3_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_wkupidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_wkupidx_1 <= io_uopin_bits_srcreq_3_wkupidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_wkupidx_1 <= s1_uop_bits_srcreq_3_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_wkupidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_wkupidx_2 <= io_uopin_bits_srcreq_3_wkupidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_wkupidx_2 <= s1_uop_bits_srcreq_3_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_wkupidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_wkupidx_3 <= io_uopin_bits_srcreq_3_wkupidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_wkupidx_3 <= s1_uop_bits_srcreq_3_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_wkupidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_wkupidx_4 <= io_uopin_bits_srcreq_3_wkupidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_wkupidx_4 <= s1_uop_bits_srcreq_3_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_3_wkupidx_5 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_3_wkupidx_5 <= io_uopin_bits_srcreq_3_wkupidx_5;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_3_wkupidx_5 <= s1_uop_bits_srcreq_3_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_valid <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_valid <= io_uopin_bits_srcreq_4_valid;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_valid <= s1_uop_bits_srcreq_4_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_isgroup <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_isgroup <= io_uopin_bits_srcreq_4_isgroup;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_iscoef <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_iscoef <= io_uopin_bits_srcreq_4_iscoef;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_idx <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_idx <= io_uopin_bits_srcreq_4_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_busy <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_busy <= io_uopin_bits_srcreq_4_busy;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_busy <= s1_uop_bits_srcreq_4_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_wkupidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_wkupidx_0 <= io_uopin_bits_srcreq_4_wkupidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_wkupidx_0 <= s1_uop_bits_srcreq_4_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_wkupidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_wkupidx_1 <= io_uopin_bits_srcreq_4_wkupidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_wkupidx_1 <= s1_uop_bits_srcreq_4_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_wkupidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_wkupidx_2 <= io_uopin_bits_srcreq_4_wkupidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_wkupidx_2 <= s1_uop_bits_srcreq_4_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_wkupidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_wkupidx_3 <= io_uopin_bits_srcreq_4_wkupidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_wkupidx_3 <= s1_uop_bits_srcreq_4_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_wkupidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_wkupidx_4 <= io_uopin_bits_srcreq_4_wkupidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_wkupidx_4 <= s1_uop_bits_srcreq_4_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_4_wkupidx_5 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_4_wkupidx_5 <= io_uopin_bits_srcreq_4_wkupidx_5;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_4_wkupidx_5 <= s1_uop_bits_srcreq_4_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_valid <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_valid <= io_uopin_bits_srcreq_5_valid;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_valid <= s1_uop_bits_srcreq_5_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_isgroup <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_isgroup <= io_uopin_bits_srcreq_5_isgroup;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_iscoef <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_iscoef <= io_uopin_bits_srcreq_5_iscoef;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_idx <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_idx <= io_uopin_bits_srcreq_5_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_busy <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_busy <= io_uopin_bits_srcreq_5_busy;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_busy <= s1_uop_bits_srcreq_5_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_wkupidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_wkupidx_0 <= io_uopin_bits_srcreq_5_wkupidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_wkupidx_0 <= s1_uop_bits_srcreq_5_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_wkupidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_wkupidx_1 <= io_uopin_bits_srcreq_5_wkupidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_wkupidx_1 <= s1_uop_bits_srcreq_5_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_wkupidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_wkupidx_2 <= io_uopin_bits_srcreq_5_wkupidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_wkupidx_2 <= s1_uop_bits_srcreq_5_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_wkupidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_wkupidx_3 <= io_uopin_bits_srcreq_5_wkupidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_wkupidx_3 <= s1_uop_bits_srcreq_5_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_wkupidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_wkupidx_4 <= io_uopin_bits_srcreq_5_wkupidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_wkupidx_4 <= s1_uop_bits_srcreq_5_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_5_wkupidx_5 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_srcreq_5_wkupidx_5 <= io_uopin_bits_srcreq_5_wkupidx_5;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_srcreq_5_wkupidx_5 <= s1_uop_bits_srcreq_5_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wbvld <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wbvld <= io_uopin_bits_wbvld;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wbreq <= 6'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wbreq <= io_uopin_bits_wbreq;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_waridx_0 <= io_uopin_bits_waridx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_waridx_0 <= out_1_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_waridx_1 <= io_uopin_bits_waridx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_waridx_1 <= out_1_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_waridx_2 <= io_uopin_bits_waridx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_waridx_2 <= out_1_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_waridx_3 <= io_uopin_bits_waridx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_waridx_3 <= out_1_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_waridx_4 <= io_uopin_bits_waridx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_waridx_4 <= out_1_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_0 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wawidx_0 <= io_uopin_bits_wawidx_0;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_wawidx_0 <= out__0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_1 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wawidx_1 <= io_uopin_bits_wawidx_1;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_wawidx_1 <= out__1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_2 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wawidx_2 <= io_uopin_bits_wawidx_2;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_wawidx_2 <= out__2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_3 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wawidx_3 <= io_uopin_bits_wawidx_3;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_wawidx_3 <= out__3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_4 <= 1'h0;
    end else if (_s1_nxt_state_T) begin
      s1_uop_bits_wawidx_4 <= io_uopin_bits_wawidx_4;
    end else if (_req2_idx_T | _T | s1_state == 2'h3) begin
      s1_uop_bits_wawidx_4 <= out__4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_state <= 2'h0;
    end else if (s1_state == 2'h0) begin
      if (_s1_nxt_state_T) begin
        if (io_uopin_bits_select | io_uopin_bits_loop) begin
          s1_state <= 2'h1;
        end else begin
          s1_state <= 2'h2;
        end
      end else begin
        s1_state <= 2'h0;
      end
    end else if (_req2_idx_T) begin
      if (read_en) begin
        s1_state <= 2'h2;
      end else begin
        s1_state <= 2'h1;
      end
    end else if (_T) begin
      if (_s1_uop_bits_srcreq_5_out_valid_T_1 & read_en) begin
        s1_state <= _s1_nxt_state_T_5;
      end
    end else if (_T_5) begin
      s1_state <= _s1_nxt_state_T_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_vld <= 1'h0;
    end else begin
      s2_vld <= read_en & s1_uop_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_wb <= 1'h0;
    end else begin
      s2_wb <= io_flop;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_wbidx <= 6'h0;
    end else begin
      s2_wbidx <= s1_uop_bits_wbreq;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_data_0 <= 32'h0;
    end else if (read_en) begin
      if (s1_uop_bits_loop & start) begin
        s2_data_0 <= loop_data;
      end else if (s1_uop_bits_drc) begin
        if (_drc_data_T_1[31]) begin
          s2_data_0 <= 32'h0;
        end else begin
          s2_data_0 <= _drc_data_T_1;
        end
      end else if (s1_uop_bits_pow) begin
        s2_data_0 <= s1_data_0_out;
      end else begin
        s2_data_0 <= io_rfreq_0_resp;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_data_1 <= 32'h0;
    end else if (read_en) begin
      if (s1_uop_bits_drcgain & ~drccoef_drcen) begin
        s2_data_1 <= 32'h800000;
      end else begin
        s2_data_1 <= io_rfreq_1_resp;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_data_2 <= 32'h0;
    end else if (start) begin
      if (s1_uop_bits_drc) begin
        if (drc1) begin
          s2_data_2 <= io_coef_mainch_drc_offset;
        end else begin
          s2_data_2 <= io_coef_subch_drc_offset;
        end
      end else begin
        s2_data_2 <= 32'h0;
      end
    end else begin
      s2_data_2 <= s2_dout;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      select <= 1'h0;
    end else if (_req2_idx_T & read_en & s1_uop_bits_select) begin
      select <= data_diff[31];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      loop_data <= 32'h0;
    end else if (_select_T_1 & s1_uop_bits_loop) begin
      if (io_coef_mainch_ch0_autoloop) begin
        loop_data <= data_diff;
      end else begin
        loop_data <= io_rfreq_0_resp;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      start <= 1'h0;
    end else begin
      start <= _s1_nxt_state_T | _GEN_214;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_uop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_uop_bits_vlen = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  s1_uop_bits_select = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_uop_bits_drc = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s1_uop_bits_pow = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s1_uop_bits_loop = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s1_uop_bits_drcgain = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s1_uop_bits_drcnum = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_isgroup = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_iscoef = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_idx = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_busy = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_3 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_4 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_5 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_isgroup = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_iscoef = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_idx = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_busy = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_valid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_isgroup = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_iscoef = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_idx = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_busy = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_wkupidx_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_wkupidx_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_wkupidx_2 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_wkupidx_3 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_wkupidx_4 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  s1_uop_bits_srcreq_2_wkupidx_5 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_isgroup = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_iscoef = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_idx = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_busy = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_wkupidx_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_wkupidx_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_wkupidx_2 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_wkupidx_3 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_wkupidx_4 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  s1_uop_bits_srcreq_3_wkupidx_5 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_valid = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_isgroup = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_iscoef = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_idx = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_busy = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_wkupidx_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_wkupidx_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_wkupidx_2 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_wkupidx_3 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_wkupidx_4 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  s1_uop_bits_srcreq_4_wkupidx_5 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_isgroup = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_iscoef = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_idx = _RAND_66[5:0];
  _RAND_67 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_busy = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_wkupidx_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_wkupidx_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_wkupidx_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_wkupidx_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_wkupidx_4 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  s1_uop_bits_srcreq_5_wkupidx_5 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  s1_uop_bits_wbvld = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  s1_uop_bits_wbreq = _RAND_75[5:0];
  _RAND_76 = {1{`RANDOM}};
  s1_uop_bits_waridx_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  s1_uop_bits_waridx_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  s1_uop_bits_waridx_2 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  s1_uop_bits_waridx_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  s1_uop_bits_waridx_4 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  s1_uop_bits_wawidx_0 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  s1_uop_bits_wawidx_1 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  s1_uop_bits_wawidx_2 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  s1_uop_bits_wawidx_3 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  s1_uop_bits_wawidx_4 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  s1_state = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  s2_vld = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  s2_wb = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  s2_wbidx = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  s2_data_0 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  s2_data_1 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  s2_data_2 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  select = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  loop_data = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  start = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  io_fwd_wkup_valid_REG = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  io_wbreq_vld_REG = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  io_wbreq_gregidx_REG = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  io_wbreq_wdata1_REG = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  io_wbreq_wdata2_REG = _RAND_100[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    s1_uop_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_vlen = 3'h0;
  end
  if (reset) begin
    s1_uop_bits_select = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_drc = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_pow = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_loop = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_drcgain = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_drcnum = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_isgroup = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_iscoef = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_isgroup = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_iscoef = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_isgroup = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_iscoef = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_2_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_isgroup = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_iscoef = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_3_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_isgroup = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_iscoef = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_4_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_isgroup = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_iscoef = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_5_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wbvld = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wbreq = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_4 = 1'h0;
  end
  if (reset) begin
    s1_state = 2'h0;
  end
  if (reset) begin
    s2_vld = 1'h0;
  end
  if (reset) begin
    s2_wb = 1'h0;
  end
  if (reset) begin
    s2_wbidx = 6'h0;
  end
  if (reset) begin
    s2_data_0 = 32'h0;
  end
  if (reset) begin
    s2_data_1 = 32'h0;
  end
  if (reset) begin
    s2_data_2 = 32'h0;
  end
  if (reset) begin
    select = 1'h0;
  end
  if (reset) begin
    loop_data = 32'h0;
  end
  if (reset) begin
    start = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Iterator(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'shc085f16) : $signed(37'sh1810be2c); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [29:0] _xtmp_T = io_din_1[36:7]; // @[coru.scala 27:26]
  wire [36:0] _GEN_0 = {{7{_xtmp_T[29]}},_xtmp_T}; // @[coru.scala 27:19]
  wire [36:0] xtmp = $signed(io_din_1) - $signed(_GEN_0); // @[coru.scala 27:19]
  wire [29:0] _ytmp_T = io_din_0[36:7]; // @[coru.scala 28:26]
  wire [36:0] _GEN_1 = {{7{_ytmp_T[29]}},_ytmp_T}; // @[coru.scala 28:19]
  wire [36:0] ytmp = $signed(io_din_0) - $signed(_GEN_1); // @[coru.scala 28:19]
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_1(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sha84de67) : $signed(37'sh1509bcce); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [30:0] _xtmp_T = io_din_1[36:6]; // @[coru.scala 27:26]
  wire [36:0] _GEN_0 = {{6{_xtmp_T[30]}},_xtmp_T}; // @[coru.scala 27:19]
  wire [36:0] xtmp = $signed(io_din_1) - $signed(_GEN_0); // @[coru.scala 27:19]
  wire [30:0] _ytmp_T = io_din_0[36:6]; // @[coru.scala 28:26]
  wire [36:0] _GEN_1 = {{6{_ytmp_T[30]}},_ytmp_T}; // @[coru.scala 28:19]
  wire [36:0] ytmp = $signed(io_din_0) - $signed(_GEN_1); // @[coru.scala 28:19]
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_2(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh8ff27e9) : $signed(37'sh11fe4fd3); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [31:0] _xtmp_T = io_din_1[36:5]; // @[coru.scala 27:26]
  wire [36:0] _GEN_0 = {{5{_xtmp_T[31]}},_xtmp_T}; // @[coru.scala 27:19]
  wire [36:0] xtmp = $signed(io_din_1) - $signed(_GEN_0); // @[coru.scala 27:19]
  wire [31:0] _ytmp_T = io_din_0[36:5]; // @[coru.scala 28:26]
  wire [36:0] _GEN_1 = {{5{_ytmp_T[31]}},_ytmp_T}; // @[coru.scala 28:19]
  wire [36:0] ytmp = $signed(io_din_0) - $signed(_GEN_1); // @[coru.scala 28:19]
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_3(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh774f166) : $signed(37'shee9e2cd); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [32:0] _xtmp_T = io_din_1[36:4]; // @[coru.scala 27:26]
  wire [36:0] _GEN_0 = {{4{_xtmp_T[32]}},_xtmp_T}; // @[coru.scala 27:19]
  wire [36:0] xtmp = $signed(io_din_1) - $signed(_GEN_0); // @[coru.scala 27:19]
  wire [32:0] _ytmp_T = io_din_0[36:4]; // @[coru.scala 28:26]
  wire [36:0] _GEN_1 = {{4{_ytmp_T[32]}},_ytmp_T}; // @[coru.scala 28:19]
  wire [36:0] ytmp = $signed(io_din_0) - $signed(_GEN_1); // @[coru.scala 28:19]
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_4(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh5e16595) : $signed(37'shbc2cb2b); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [33:0] _xtmp_T = io_din_1[36:3]; // @[coru.scala 27:26]
  wire [36:0] _GEN_0 = {{3{_xtmp_T[33]}},_xtmp_T}; // @[coru.scala 27:19]
  wire [36:0] xtmp = $signed(io_din_1) - $signed(_GEN_0); // @[coru.scala 27:19]
  wire [33:0] _ytmp_T = io_din_0[36:3]; // @[coru.scala 28:26]
  wire [36:0] _GEN_1 = {{3{_ytmp_T[33]}},_ytmp_T}; // @[coru.scala 28:19]
  wire [36:0] ytmp = $signed(io_din_0) - $signed(_GEN_1); // @[coru.scala 28:19]
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_5(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh439b9ba) : $signed(37'sh8737374); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [34:0] _xtmp_T = io_din_1[36:2]; // @[coru.scala 27:26]
  wire [36:0] _GEN_0 = {{2{_xtmp_T[34]}},_xtmp_T}; // @[coru.scala 27:19]
  wire [36:0] xtmp = $signed(io_din_1) - $signed(_GEN_0); // @[coru.scala 27:19]
  wire [34:0] _ytmp_T = io_din_0[36:2]; // @[coru.scala 28:26]
  wire [36:0] _GEN_1 = {{2{_ytmp_T[34]}},_ytmp_T}; // @[coru.scala 28:19]
  wire [36:0] ytmp = $signed(io_din_0) - $signed(_GEN_1); // @[coru.scala 28:19]
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_6(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh262b718) : $signed(37'sh4c56e2f); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [35:0] _xtmp_T = io_din_1[36:1]; // @[coru.scala 24:20]
  wire [35:0] _ytmp_T = io_din_0[36:1]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{1{_xtmp_T[35]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{1{_ytmp_T[35]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_7(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh11bf766) : $signed(37'sh237eecc); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [34:0] _xtmp_T = io_din_1[36:2]; // @[coru.scala 24:20]
  wire [34:0] _ytmp_T = io_din_0[36:2]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{2{_xtmp_T[34]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{2{_ytmp_T[34]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_8(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh8bb476) : $signed(37'sh11768eb); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [33:0] _xtmp_T = io_din_1[36:3]; // @[coru.scala 24:20]
  wire [33:0] _ytmp_T = io_din_0[36:3]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{3{_xtmp_T[33]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{3{_ytmp_T[33]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_9(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh4593eb) : $signed(37'sh8b27d6); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [32:0] _xtmp_T = io_din_1[36:4]; // @[coru.scala 24:20]
  wire [32:0] _ytmp_T = io_din_0[36:4]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{4{_xtmp_T[32]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{4{_ytmp_T[32]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_11(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh22c13f) : $signed(37'sh45827f); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [31:0] _xtmp_T = io_din_1[36:5]; // @[coru.scala 24:20]
  wire [31:0] _ytmp_T = io_din_0[36:5]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{5{_xtmp_T[31]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{5{_ytmp_T[31]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_12(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh115f8a) : $signed(37'sh22bf13); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [30:0] _xtmp_T = io_din_1[36:6]; // @[coru.scala 24:20]
  wire [30:0] _ytmp_T = io_din_0[36:6]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{6{_xtmp_T[30]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{6{_ytmp_T[30]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_13(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh8afa2) : $signed(37'sh115f44); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [29:0] _xtmp_T = io_din_1[36:7]; // @[coru.scala 24:20]
  wire [29:0] _ytmp_T = io_din_0[36:7]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{7{_xtmp_T[29]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{7{_ytmp_T[29]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_14(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_1,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh457cd) : $signed(37'sh8af99); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [28:0] _xtmp_T = io_din_1[36:8]; // @[coru.scala 24:20]
  wire [28:0] _ytmp_T = io_din_0[36:8]; // @[coru.scala 25:20]
  wire [36:0] xtmp = {{8{_xtmp_T[28]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] ytmp = {{8{_ytmp_T[28]}},_ytmp_T};
  wire [36:0] _yout_T_2 = $signed(io_din_1) + $signed(ytmp); // @[coru.scala 32:29]
  wire [36:0] _yout_T_5 = $signed(io_din_1) - $signed(ytmp); // @[coru.scala 32:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_1 = sel ? $signed(_yout_T_2) : $signed(_yout_T_5); // @[coru.scala 32:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module Iterator_15(
  input  [36:0] io_din_0,
  input  [36:0] io_din_1,
  input  [36:0] io_din_2,
  output [36:0] io_dout_0,
  output [36:0] io_dout_2,
  input         io_cortype
);
  wire [36:0] dzin = io_cortype ? $signed(37'sh22be6) : $signed(37'sh457cc); // @[coru.scala 38:17]
  wire  sel = io_cortype ? ~io_din_2[36] : io_din_1[36]; // @[coru.scala 39:17]
  wire [27:0] _xtmp_T = io_din_1[36:9]; // @[coru.scala 24:20]
  wire [36:0] xtmp = {{9{_xtmp_T[27]}},_xtmp_T};
  wire [36:0] _xout_T_2 = $signed(io_din_0) + $signed(xtmp); // @[coru.scala 31:29]
  wire [36:0] _xout_T_5 = $signed(io_din_0) - $signed(xtmp); // @[coru.scala 31:41]
  wire [36:0] _zout_T_2 = $signed(io_din_2) - $signed(dzin); // @[coru.scala 33:29]
  wire [36:0] _zout_T_5 = $signed(io_din_2) + $signed(dzin); // @[coru.scala 33:41]
  assign io_dout_0 = sel ? $signed(_xout_T_2) : $signed(_xout_T_5); // @[coru.scala 31:16]
  assign io_dout_2 = sel ? $signed(_zout_T_2) : $signed(_zout_T_5); // @[coru.scala 33:16]
endmodule
module CorUnit(
  input         clock,
  input         reset,
  output        io_uopin_ready,
  input         io_uopin_valid,
  input         io_uopin_bits_cortype,
  input         io_uopin_bits_srcreq_0_valid,
  input  [5:0]  io_uopin_bits_srcreq_0_idx,
  input         io_uopin_bits_srcreq_0_busy,
  input         io_uopin_bits_srcreq_0_wkupidx_0,
  input         io_uopin_bits_srcreq_0_wkupidx_1,
  input         io_uopin_bits_srcreq_0_wkupidx_2,
  input         io_uopin_bits_srcreq_0_wkupidx_3,
  input         io_uopin_bits_srcreq_0_wkupidx_4,
  input         io_uopin_bits_srcreq_0_wkupidx_5,
  input         io_uopin_bits_srcreq_1_valid,
  input  [5:0]  io_uopin_bits_srcreq_1_idx,
  input         io_uopin_bits_srcreq_1_busy,
  input         io_uopin_bits_srcreq_1_wkupidx_0,
  input         io_uopin_bits_srcreq_1_wkupidx_1,
  input         io_uopin_bits_srcreq_1_wkupidx_2,
  input         io_uopin_bits_srcreq_1_wkupidx_3,
  input         io_uopin_bits_srcreq_1_wkupidx_4,
  input         io_uopin_bits_srcreq_1_wkupidx_5,
  input         io_uopin_bits_wbvld,
  input  [5:0]  io_uopin_bits_wbreq,
  input         io_uopin_bits_waridx_0,
  input         io_uopin_bits_waridx_1,
  input         io_uopin_bits_waridx_2,
  input         io_uopin_bits_waridx_3,
  input         io_uopin_bits_waridx_4,
  input         io_uopin_bits_wawidx_0,
  input         io_uopin_bits_wawidx_1,
  input         io_uopin_bits_wawidx_2,
  input         io_uopin_bits_wawidx_3,
  input         io_uopin_bits_wawidx_4,
  output [5:0]  io_rfreq_0_req_idx,
  input  [31:0] io_rfreq_0_resp,
  output [5:0]  io_rfreq_1_req_idx,
  input  [31:0] io_rfreq_1_resp,
  output [31:0] io_wbreq_wdata2,
  output        io_wbreq_vld,
  output [5:0]  io_wbreq_gregidx,
  output        io_empty,
  output        io_fwd_wkup_valid,
  output [5:0]  io_fwd_wkup_bits,
  input         io_raw_wkup_0_valid,
  input  [5:0]  io_raw_wkup_0_bits,
  input         io_raw_wkup_1_valid,
  input  [5:0]  io_raw_wkup_1_bits,
  input         io_raw_wkup_2_valid,
  input  [5:0]  io_raw_wkup_2_bits,
  input         io_raw_wkup_3_valid,
  input  [5:0]  io_raw_wkup_3_bits,
  input         io_raw_wkup_4_valid,
  input  [5:0]  io_raw_wkup_4_bits,
  input         io_raw_wkup_5_valid,
  input  [5:0]  io_raw_wkup_5_bits,
  output        io_wbcheck_valid,
  output [5:0]  io_wbcheck_bits,
  output        io_r_check_0_valid,
  output [5:0]  io_r_check_0_bits,
  output        io_r_check_1_valid,
  output [5:0]  io_r_check_1_bits,
  input         io_other_flop_0,
  input         io_other_flop_1,
  input         io_other_flop_2,
  input         io_other_flop_3,
  input         io_other_flop_4,
  output        io_flop
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire [36:0] inst_io_din_0; // @[coru.scala 165:22]
  wire [36:0] inst_io_din_1; // @[coru.scala 165:22]
  wire [36:0] inst_io_din_2; // @[coru.scala 165:22]
  wire [36:0] inst_io_dout_0; // @[coru.scala 165:22]
  wire [36:0] inst_io_dout_1; // @[coru.scala 165:22]
  wire [36:0] inst_io_dout_2; // @[coru.scala 165:22]
  wire  inst_io_cortype; // @[coru.scala 165:22]
  wire [36:0] inst_1_io_din_0; // @[coru.scala 165:22]
  wire [36:0] inst_1_io_din_1; // @[coru.scala 165:22]
  wire [36:0] inst_1_io_din_2; // @[coru.scala 165:22]
  wire [36:0] inst_1_io_dout_0; // @[coru.scala 165:22]
  wire [36:0] inst_1_io_dout_1; // @[coru.scala 165:22]
  wire [36:0] inst_1_io_dout_2; // @[coru.scala 165:22]
  wire  inst_1_io_cortype; // @[coru.scala 165:22]
  wire [36:0] inst_2_io_din_0; // @[coru.scala 165:22]
  wire [36:0] inst_2_io_din_1; // @[coru.scala 165:22]
  wire [36:0] inst_2_io_din_2; // @[coru.scala 165:22]
  wire [36:0] inst_2_io_dout_0; // @[coru.scala 165:22]
  wire [36:0] inst_2_io_dout_1; // @[coru.scala 165:22]
  wire [36:0] inst_2_io_dout_2; // @[coru.scala 165:22]
  wire  inst_2_io_cortype; // @[coru.scala 165:22]
  wire [36:0] inst_3_io_din_0; // @[coru.scala 165:22]
  wire [36:0] inst_3_io_din_1; // @[coru.scala 165:22]
  wire [36:0] inst_3_io_din_2; // @[coru.scala 165:22]
  wire [36:0] inst_3_io_dout_0; // @[coru.scala 165:22]
  wire [36:0] inst_3_io_dout_1; // @[coru.scala 165:22]
  wire [36:0] inst_3_io_dout_2; // @[coru.scala 165:22]
  wire  inst_3_io_cortype; // @[coru.scala 165:22]
  wire [36:0] inst_4_io_din_0; // @[coru.scala 165:22]
  wire [36:0] inst_4_io_din_1; // @[coru.scala 165:22]
  wire [36:0] inst_4_io_din_2; // @[coru.scala 165:22]
  wire [36:0] inst_4_io_dout_0; // @[coru.scala 165:22]
  wire [36:0] inst_4_io_dout_1; // @[coru.scala 165:22]
  wire [36:0] inst_4_io_dout_2; // @[coru.scala 165:22]
  wire  inst_4_io_cortype; // @[coru.scala 165:22]
  wire [36:0] inst_5_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_5_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_5_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_5_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_5_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_5_io_dout_2; // @[coru.scala 199:22]
  wire  inst_5_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_6_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_6_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_6_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_6_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_6_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_6_io_dout_2; // @[coru.scala 199:22]
  wire  inst_6_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_7_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_7_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_7_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_7_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_7_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_7_io_dout_2; // @[coru.scala 199:22]
  wire  inst_7_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_8_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_8_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_8_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_8_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_8_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_8_io_dout_2; // @[coru.scala 199:22]
  wire  inst_8_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_9_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_9_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_9_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_9_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_9_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_9_io_dout_2; // @[coru.scala 199:22]
  wire  inst_9_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_10_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_10_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_10_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_10_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_10_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_10_io_dout_2; // @[coru.scala 199:22]
  wire  inst_10_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_11_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_11_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_11_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_11_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_11_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_11_io_dout_2; // @[coru.scala 199:22]
  wire  inst_11_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_12_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_12_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_12_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_12_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_12_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_12_io_dout_2; // @[coru.scala 199:22]
  wire  inst_12_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_13_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_13_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_13_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_13_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_13_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_13_io_dout_2; // @[coru.scala 199:22]
  wire  inst_13_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_14_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_14_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_14_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_14_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_14_io_dout_1; // @[coru.scala 199:22]
  wire [36:0] inst_14_io_dout_2; // @[coru.scala 199:22]
  wire  inst_14_io_cortype; // @[coru.scala 199:22]
  wire [36:0] inst_15_io_din_0; // @[coru.scala 199:22]
  wire [36:0] inst_15_io_din_1; // @[coru.scala 199:22]
  wire [36:0] inst_15_io_din_2; // @[coru.scala 199:22]
  wire [36:0] inst_15_io_dout_0; // @[coru.scala 199:22]
  wire [36:0] inst_15_io_dout_2; // @[coru.scala 199:22]
  wire  inst_15_io_cortype; // @[coru.scala 199:22]
  reg  s1_uop_valid; // @[coru.scala 64:24]
  reg  s1_uop_bits_cortype; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_valid; // @[coru.scala 64:24]
  reg [5:0] s1_uop_bits_srcreq_0_idx; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_busy; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_wkupidx_0; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_wkupidx_1; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_wkupidx_2; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_wkupidx_3; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_wkupidx_4; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_0_wkupidx_5; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_valid; // @[coru.scala 64:24]
  reg [5:0] s1_uop_bits_srcreq_1_idx; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_busy; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_wkupidx_0; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_wkupidx_1; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_wkupidx_2; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_wkupidx_3; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_wkupidx_4; // @[coru.scala 64:24]
  reg  s1_uop_bits_srcreq_1_wkupidx_5; // @[coru.scala 64:24]
  reg  s1_uop_bits_wbvld; // @[coru.scala 64:24]
  reg [5:0] s1_uop_bits_wbreq; // @[coru.scala 64:24]
  reg  s1_uop_bits_waridx_0; // @[coru.scala 64:24]
  reg  s1_uop_bits_waridx_1; // @[coru.scala 64:24]
  reg  s1_uop_bits_waridx_2; // @[coru.scala 64:24]
  reg  s1_uop_bits_waridx_3; // @[coru.scala 64:24]
  reg  s1_uop_bits_waridx_4; // @[coru.scala 64:24]
  reg  s1_uop_bits_wawidx_0; // @[coru.scala 64:24]
  reg  s1_uop_bits_wawidx_1; // @[coru.scala 64:24]
  reg  s1_uop_bits_wawidx_2; // @[coru.scala 64:24]
  reg  s1_uop_bits_wawidx_3; // @[coru.scala 64:24]
  reg  s1_uop_bits_wawidx_4; // @[coru.scala 64:24]
  reg  s2_vld; // @[coru.scala 65:24]
  reg [5:0] s2_wbidx; // @[coru.scala 66:25]
  wire  _no_depd_T_7 = s1_uop_bits_wawidx_0 | s1_uop_bits_wawidx_1 | s1_uop_bits_wawidx_2 | s1_uop_bits_wawidx_3 |
    s1_uop_bits_wawidx_4; // @[coru.scala 68:46]
  wire  no_depd = ~(s1_uop_bits_waridx_0 | s1_uop_bits_waridx_1 | s1_uop_bits_waridx_2 | s1_uop_bits_waridx_3 |
    s1_uop_bits_waridx_4 | _no_depd_T_7); // @[coru.scala 67:17]
  wire  read_en = (s1_uop_bits_srcreq_0_valid & ~s1_uop_bits_srcreq_0_busy | ~s1_uop_bits_srcreq_0_valid) & (
    s1_uop_bits_srcreq_1_valid & ~s1_uop_bits_srcreq_1_busy | ~s1_uop_bits_srcreq_1_valid); // @[coru.scala 135:82]
  wire  flop = no_depd & read_en & s1_uop_valid; // @[coru.scala 117:33]
  wire  s1_uop_bits_srcreq_0_out_valid = s1_uop_bits_srcreq_0_valid & ~io_flop; // @[coru.scala 73:28]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_0_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_0_out_wkupidx_0_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_0 = s1_uop_bits_srcreq_0_wkupidx_0 & _s1_uop_bits_srcreq_0_out_wkupidx_0_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_0_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_0_out_wkupidx_1_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_1 = s1_uop_bits_srcreq_0_wkupidx_1 & _s1_uop_bits_srcreq_0_out_wkupidx_1_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_0_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_0_out_wkupidx_2_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_2 = s1_uop_bits_srcreq_0_wkupidx_2 & _s1_uop_bits_srcreq_0_out_wkupidx_2_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_0_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_0_out_wkupidx_3_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_3 = s1_uop_bits_srcreq_0_wkupidx_3 & _s1_uop_bits_srcreq_0_out_wkupidx_3_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_0_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_0_out_wkupidx_4_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_4 = s1_uop_bits_srcreq_0_wkupidx_4 & _s1_uop_bits_srcreq_0_out_wkupidx_4_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_0_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_0_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_0_out_wkupidx_5_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_0_out_wkupidx_5 = s1_uop_bits_srcreq_0_wkupidx_5 & _s1_uop_bits_srcreq_0_out_wkupidx_5_T_2; // @[coru.scala 75:40]
  wire  s1_uop_bits_srcreq_0_out_busy = s1_uop_bits_srcreq_0_out_wkupidx_0 | s1_uop_bits_srcreq_0_out_wkupidx_1 |
    s1_uop_bits_srcreq_0_out_wkupidx_2 | s1_uop_bits_srcreq_0_out_wkupidx_3 | s1_uop_bits_srcreq_0_out_wkupidx_4 |
    s1_uop_bits_srcreq_0_out_wkupidx_5; // @[coru.scala 79:37]
  wire  s1_uop_bits_srcreq_1_out_valid = s1_uop_bits_srcreq_1_valid & ~io_flop; // @[coru.scala 73:28]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_0_T_1 = io_raw_wkup_0_bits != s1_uop_bits_srcreq_1_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_0_T_2 = ~io_raw_wkup_0_valid | _s1_uop_bits_srcreq_1_out_wkupidx_0_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_0 = s1_uop_bits_srcreq_1_wkupidx_0 & _s1_uop_bits_srcreq_1_out_wkupidx_0_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_1_T_1 = io_raw_wkup_1_bits != s1_uop_bits_srcreq_1_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_1_T_2 = ~io_raw_wkup_1_valid | _s1_uop_bits_srcreq_1_out_wkupidx_1_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_1 = s1_uop_bits_srcreq_1_wkupidx_1 & _s1_uop_bits_srcreq_1_out_wkupidx_1_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_2_T_1 = io_raw_wkup_2_bits != s1_uop_bits_srcreq_1_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_2_T_2 = ~io_raw_wkup_2_valid | _s1_uop_bits_srcreq_1_out_wkupidx_2_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_2 = s1_uop_bits_srcreq_1_wkupidx_2 & _s1_uop_bits_srcreq_1_out_wkupidx_2_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_3_T_1 = io_raw_wkup_3_bits != s1_uop_bits_srcreq_1_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_3_T_2 = ~io_raw_wkup_3_valid | _s1_uop_bits_srcreq_1_out_wkupidx_3_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_3 = s1_uop_bits_srcreq_1_wkupidx_3 & _s1_uop_bits_srcreq_1_out_wkupidx_3_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_4_T_1 = io_raw_wkup_4_bits != s1_uop_bits_srcreq_1_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_4_T_2 = ~io_raw_wkup_4_valid | _s1_uop_bits_srcreq_1_out_wkupidx_4_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_4 = s1_uop_bits_srcreq_1_wkupidx_4 & _s1_uop_bits_srcreq_1_out_wkupidx_4_T_2; // @[coru.scala 75:40]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_5_T_1 = io_raw_wkup_5_bits != s1_uop_bits_srcreq_1_idx; // @[coru.scala 77:32]
  wire  _s1_uop_bits_srcreq_1_out_wkupidx_5_T_2 = ~io_raw_wkup_5_valid | _s1_uop_bits_srcreq_1_out_wkupidx_5_T_1; // @[coru.scala 76:32]
  wire  s1_uop_bits_srcreq_1_out_wkupidx_5 = s1_uop_bits_srcreq_1_wkupidx_5 & _s1_uop_bits_srcreq_1_out_wkupidx_5_T_2; // @[coru.scala 75:40]
  wire  s1_uop_bits_srcreq_1_out_busy = s1_uop_bits_srcreq_1_out_wkupidx_0 | s1_uop_bits_srcreq_1_out_wkupidx_1 |
    s1_uop_bits_srcreq_1_out_wkupidx_2 | s1_uop_bits_srcreq_1_out_wkupidx_3 | s1_uop_bits_srcreq_1_out_wkupidx_4 |
    s1_uop_bits_srcreq_1_out_wkupidx_5; // @[coru.scala 79:37]
  wire  out__0 = s1_uop_bits_waridx_0 & ~io_other_flop_0; // @[coru.scala 85:41]
  wire  out__1 = s1_uop_bits_waridx_1 & ~io_other_flop_1; // @[coru.scala 85:41]
  wire  out__2 = s1_uop_bits_waridx_2 & ~io_other_flop_2; // @[coru.scala 85:41]
  wire  out__3 = s1_uop_bits_waridx_3 & ~io_other_flop_3; // @[coru.scala 85:41]
  wire  out__4 = s1_uop_bits_waridx_4 & ~io_other_flop_4; // @[coru.scala 85:41]
  wire  out_1_0 = s1_uop_bits_wawidx_0 & ~io_other_flop_0; // @[coru.scala 85:41]
  wire  out_1_1 = s1_uop_bits_wawidx_1 & ~io_other_flop_1; // @[coru.scala 85:41]
  wire  out_1_2 = s1_uop_bits_wawidx_2 & ~io_other_flop_2; // @[coru.scala 85:41]
  wire  out_1_3 = s1_uop_bits_wawidx_3 & ~io_other_flop_3; // @[coru.scala 85:41]
  wire  out_1_4 = s1_uop_bits_wawidx_4 & ~io_other_flop_4; // @[coru.scala 85:41]
  wire  _io_wbcheck_valid_T = ~flop; // @[coru.scala 138:39]
  wire  _io_empty_T = ~s1_uop_valid; // @[coru.scala 147:15]
  wire [31:0] _T_20 = io_rfreq_0_resp; // @[coru.scala 153:47]
  wire [31:0] _T_21 = io_rfreq_1_resp; // @[coru.scala 153:47]
  wire [36:0] rf_resp_0 = {{5{_T_20[31]}},_T_20}; // @[coru.scala 153:47 coru.scala 153:47]
  wire [36:0] rf_resp_1 = {{5{_T_21[31]}},_T_21}; // @[coru.scala 153:47 coru.scala 153:47]
  wire [36:0] _maxdata_T_2 = $signed(rf_resp_0) - $signed(rf_resp_1); // @[coru.scala 155:33]
  wire [36:0] maxdata = _maxdata_T_2[36] ? $signed(rf_resp_1) : $signed(rf_resp_0); // @[coru.scala 155:20]
  wire [36:0] _s1_data_0_0_T_2 = $signed(maxdata) + 37'sh800000; // @[coru.scala 159:66]
  wire [36:0] _s1_data_0_1_T_2 = $signed(maxdata) - 37'sh800000; // @[coru.scala 160:66]
  wire  _T_22 = io_uopin_ready & io_uopin_valid; // @[Decoupled.scala 40:37]
  wire  _s2_vld_T = s1_uop_valid & flop; // @[coru.scala 183:26]
  reg  s2_cortype; // @[coru.scala 190:27]
  reg [36:0] s1_data_reg_0; // @[coru.scala 191:28]
  reg [36:0] s1_data_reg_1; // @[coru.scala 191:28]
  reg [36:0] s1_data_reg_2; // @[coru.scala 191:28]
  wire [36:0] s1_data_5_0 = inst_4_io_dout_0; // @[coru.scala 151:24 coru.scala 167:18]
  wire [36:0] s1_data_5_1 = inst_4_io_dout_1; // @[coru.scala 151:24 coru.scala 167:18]
  wire [36:0] s1_data_5_2 = inst_4_io_dout_2; // @[coru.scala 151:24 coru.scala 167:18]
  wire [36:0] s2_data_11_0 = inst_15_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  wire [36:0] s2_data_11_2 = inst_15_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  wire [36:0] s2_out = s2_cortype ? $signed(s2_data_11_0) : $signed(s2_data_11_2); // @[coru.scala 206:19]
  reg  io_wbreq_vld_REG; // @[coru.scala 211:26]
  reg [5:0] io_wbreq_gregidx_REG; // @[coru.scala 212:30]
  reg [31:0] io_wbreq_wdata2_REG; // @[coru.scala 214:29]
  Iterator inst ( // @[coru.scala 165:22]
    .io_din_0(inst_io_din_0),
    .io_din_1(inst_io_din_1),
    .io_din_2(inst_io_din_2),
    .io_dout_0(inst_io_dout_0),
    .io_dout_1(inst_io_dout_1),
    .io_dout_2(inst_io_dout_2),
    .io_cortype(inst_io_cortype)
  );
  Iterator_1 inst_1 ( // @[coru.scala 165:22]
    .io_din_0(inst_1_io_din_0),
    .io_din_1(inst_1_io_din_1),
    .io_din_2(inst_1_io_din_2),
    .io_dout_0(inst_1_io_dout_0),
    .io_dout_1(inst_1_io_dout_1),
    .io_dout_2(inst_1_io_dout_2),
    .io_cortype(inst_1_io_cortype)
  );
  Iterator_2 inst_2 ( // @[coru.scala 165:22]
    .io_din_0(inst_2_io_din_0),
    .io_din_1(inst_2_io_din_1),
    .io_din_2(inst_2_io_din_2),
    .io_dout_0(inst_2_io_dout_0),
    .io_dout_1(inst_2_io_dout_1),
    .io_dout_2(inst_2_io_dout_2),
    .io_cortype(inst_2_io_cortype)
  );
  Iterator_3 inst_3 ( // @[coru.scala 165:22]
    .io_din_0(inst_3_io_din_0),
    .io_din_1(inst_3_io_din_1),
    .io_din_2(inst_3_io_din_2),
    .io_dout_0(inst_3_io_dout_0),
    .io_dout_1(inst_3_io_dout_1),
    .io_dout_2(inst_3_io_dout_2),
    .io_cortype(inst_3_io_cortype)
  );
  Iterator_4 inst_4 ( // @[coru.scala 165:22]
    .io_din_0(inst_4_io_din_0),
    .io_din_1(inst_4_io_din_1),
    .io_din_2(inst_4_io_din_2),
    .io_dout_0(inst_4_io_dout_0),
    .io_dout_1(inst_4_io_dout_1),
    .io_dout_2(inst_4_io_dout_2),
    .io_cortype(inst_4_io_cortype)
  );
  Iterator_5 inst_5 ( // @[coru.scala 199:22]
    .io_din_0(inst_5_io_din_0),
    .io_din_1(inst_5_io_din_1),
    .io_din_2(inst_5_io_din_2),
    .io_dout_0(inst_5_io_dout_0),
    .io_dout_1(inst_5_io_dout_1),
    .io_dout_2(inst_5_io_dout_2),
    .io_cortype(inst_5_io_cortype)
  );
  Iterator_6 inst_6 ( // @[coru.scala 199:22]
    .io_din_0(inst_6_io_din_0),
    .io_din_1(inst_6_io_din_1),
    .io_din_2(inst_6_io_din_2),
    .io_dout_0(inst_6_io_dout_0),
    .io_dout_1(inst_6_io_dout_1),
    .io_dout_2(inst_6_io_dout_2),
    .io_cortype(inst_6_io_cortype)
  );
  Iterator_7 inst_7 ( // @[coru.scala 199:22]
    .io_din_0(inst_7_io_din_0),
    .io_din_1(inst_7_io_din_1),
    .io_din_2(inst_7_io_din_2),
    .io_dout_0(inst_7_io_dout_0),
    .io_dout_1(inst_7_io_dout_1),
    .io_dout_2(inst_7_io_dout_2),
    .io_cortype(inst_7_io_cortype)
  );
  Iterator_8 inst_8 ( // @[coru.scala 199:22]
    .io_din_0(inst_8_io_din_0),
    .io_din_1(inst_8_io_din_1),
    .io_din_2(inst_8_io_din_2),
    .io_dout_0(inst_8_io_dout_0),
    .io_dout_1(inst_8_io_dout_1),
    .io_dout_2(inst_8_io_dout_2),
    .io_cortype(inst_8_io_cortype)
  );
  Iterator_9 inst_9 ( // @[coru.scala 199:22]
    .io_din_0(inst_9_io_din_0),
    .io_din_1(inst_9_io_din_1),
    .io_din_2(inst_9_io_din_2),
    .io_dout_0(inst_9_io_dout_0),
    .io_dout_1(inst_9_io_dout_1),
    .io_dout_2(inst_9_io_dout_2),
    .io_cortype(inst_9_io_cortype)
  );
  Iterator_9 inst_10 ( // @[coru.scala 199:22]
    .io_din_0(inst_10_io_din_0),
    .io_din_1(inst_10_io_din_1),
    .io_din_2(inst_10_io_din_2),
    .io_dout_0(inst_10_io_dout_0),
    .io_dout_1(inst_10_io_dout_1),
    .io_dout_2(inst_10_io_dout_2),
    .io_cortype(inst_10_io_cortype)
  );
  Iterator_11 inst_11 ( // @[coru.scala 199:22]
    .io_din_0(inst_11_io_din_0),
    .io_din_1(inst_11_io_din_1),
    .io_din_2(inst_11_io_din_2),
    .io_dout_0(inst_11_io_dout_0),
    .io_dout_1(inst_11_io_dout_1),
    .io_dout_2(inst_11_io_dout_2),
    .io_cortype(inst_11_io_cortype)
  );
  Iterator_12 inst_12 ( // @[coru.scala 199:22]
    .io_din_0(inst_12_io_din_0),
    .io_din_1(inst_12_io_din_1),
    .io_din_2(inst_12_io_din_2),
    .io_dout_0(inst_12_io_dout_0),
    .io_dout_1(inst_12_io_dout_1),
    .io_dout_2(inst_12_io_dout_2),
    .io_cortype(inst_12_io_cortype)
  );
  Iterator_13 inst_13 ( // @[coru.scala 199:22]
    .io_din_0(inst_13_io_din_0),
    .io_din_1(inst_13_io_din_1),
    .io_din_2(inst_13_io_din_2),
    .io_dout_0(inst_13_io_dout_0),
    .io_dout_1(inst_13_io_dout_1),
    .io_dout_2(inst_13_io_dout_2),
    .io_cortype(inst_13_io_cortype)
  );
  Iterator_14 inst_14 ( // @[coru.scala 199:22]
    .io_din_0(inst_14_io_din_0),
    .io_din_1(inst_14_io_din_1),
    .io_din_2(inst_14_io_din_2),
    .io_dout_0(inst_14_io_dout_0),
    .io_dout_1(inst_14_io_dout_1),
    .io_dout_2(inst_14_io_dout_2),
    .io_cortype(inst_14_io_cortype)
  );
  Iterator_15 inst_15 ( // @[coru.scala 199:22]
    .io_din_0(inst_15_io_din_0),
    .io_din_1(inst_15_io_din_1),
    .io_din_2(inst_15_io_din_2),
    .io_dout_0(inst_15_io_dout_0),
    .io_dout_2(inst_15_io_dout_2),
    .io_cortype(inst_15_io_cortype)
  );
  assign io_uopin_ready = flop | _io_empty_T; // @[coru.scala 148:26]
  assign io_rfreq_0_req_idx = s1_uop_bits_srcreq_0_idx; // @[coru.scala 130:29]
  assign io_rfreq_1_req_idx = s1_uop_bits_srcreq_1_idx; // @[coru.scala 130:29]
  assign io_wbreq_wdata2 = io_wbreq_wdata2_REG; // @[coru.scala 214:19]
  assign io_wbreq_vld = io_wbreq_vld_REG; // @[coru.scala 211:16]
  assign io_wbreq_gregidx = io_wbreq_gregidx_REG; // @[coru.scala 212:20]
  assign io_empty = ~s1_uop_valid & ~s2_vld & ~io_wbreq_vld; // @[coru.scala 147:40]
  assign io_fwd_wkup_valid = s2_vld; // @[coru.scala 186:21]
  assign io_fwd_wkup_bits = s2_wbidx; // @[coru.scala 187:20]
  assign io_wbcheck_valid = s1_uop_valid & ~flop & s1_uop_bits_wbvld; // @[coru.scala 138:45]
  assign io_wbcheck_bits = s1_uop_bits_wbreq; // @[coru.scala 139:20]
  assign io_r_check_0_valid = s1_uop_valid & s1_uop_bits_srcreq_0_valid & _io_wbcheck_valid_T; // @[coru.scala 143:54]
  assign io_r_check_0_bits = s1_uop_bits_srcreq_0_idx; // @[coru.scala 144:25]
  assign io_r_check_1_valid = s1_uop_valid & s1_uop_bits_srcreq_1_valid & _io_wbcheck_valid_T; // @[coru.scala 143:54]
  assign io_r_check_1_bits = s1_uop_bits_srcreq_1_idx; // @[coru.scala 144:25]
  assign io_flop = no_depd & read_en & s1_uop_valid; // @[coru.scala 117:33]
  assign inst_io_din_0 = s1_uop_bits_cortype ? $signed(37'sh3e25edc5f) : $signed(_s1_data_0_0_T_2); // @[coru.scala 159:23]
  assign inst_io_din_1 = s1_uop_bits_cortype ? $signed(37'sh3e25edc5f) : $signed(_s1_data_0_1_T_2); // @[coru.scala 160:23]
  assign inst_io_din_2 = s1_uop_bits_cortype ? $signed(rf_resp_0) : $signed(37'sh0); // @[coru.scala 161:23]
  assign inst_io_cortype = s1_uop_bits_cortype; // @[coru.scala 168:21]
  assign inst_1_io_din_0 = inst_io_dout_0; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_1_io_din_1 = inst_io_dout_1; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_1_io_din_2 = inst_io_dout_2; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_1_io_cortype = s1_uop_bits_cortype; // @[coru.scala 168:21]
  assign inst_2_io_din_0 = inst_1_io_dout_0; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_2_io_din_1 = inst_1_io_dout_1; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_2_io_din_2 = inst_1_io_dout_2; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_2_io_cortype = s1_uop_bits_cortype; // @[coru.scala 168:21]
  assign inst_3_io_din_0 = inst_2_io_dout_0; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_3_io_din_1 = inst_2_io_dout_1; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_3_io_din_2 = inst_2_io_dout_2; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_3_io_cortype = s1_uop_bits_cortype; // @[coru.scala 168:21]
  assign inst_4_io_din_0 = inst_3_io_dout_0; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_4_io_din_1 = inst_3_io_dout_1; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_4_io_din_2 = inst_3_io_dout_2; // @[coru.scala 151:24 coru.scala 167:18]
  assign inst_4_io_cortype = s1_uop_bits_cortype; // @[coru.scala 168:21]
  assign inst_5_io_din_0 = s1_data_reg_0; // @[coru.scala 189:24 coru.scala 193:14]
  assign inst_5_io_din_1 = s1_data_reg_1; // @[coru.scala 189:24 coru.scala 193:14]
  assign inst_5_io_din_2 = s1_data_reg_2; // @[coru.scala 189:24 coru.scala 193:14]
  assign inst_5_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_6_io_din_0 = inst_5_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_6_io_din_1 = inst_5_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_6_io_din_2 = inst_5_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_6_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_7_io_din_0 = inst_6_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_7_io_din_1 = inst_6_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_7_io_din_2 = inst_6_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_7_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_8_io_din_0 = inst_7_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_8_io_din_1 = inst_7_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_8_io_din_2 = inst_7_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_8_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_9_io_din_0 = inst_8_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_9_io_din_1 = inst_8_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_9_io_din_2 = inst_8_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_9_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_10_io_din_0 = inst_9_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_10_io_din_1 = inst_9_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_10_io_din_2 = inst_9_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_10_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_11_io_din_0 = inst_10_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_11_io_din_1 = inst_10_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_11_io_din_2 = inst_10_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_11_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_12_io_din_0 = inst_11_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_12_io_din_1 = inst_11_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_12_io_din_2 = inst_11_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_12_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_13_io_din_0 = inst_12_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_13_io_din_1 = inst_12_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_13_io_din_2 = inst_12_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_13_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_14_io_din_0 = inst_13_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_14_io_din_1 = inst_13_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_14_io_din_2 = inst_13_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_14_io_cortype = s2_cortype; // @[coru.scala 203:21]
  assign inst_15_io_din_0 = inst_14_io_dout_0; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_15_io_din_1 = inst_14_io_dout_1; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_15_io_din_2 = inst_14_io_dout_2; // @[coru.scala 189:24 coru.scala 200:18]
  assign inst_15_io_cortype = s2_cortype; // @[coru.scala 203:21]
  always @(posedge clock) begin
    io_wbreq_vld_REG <= s2_vld; // @[coru.scala 211:26]
    io_wbreq_gregidx_REG <= s2_wbidx; // @[coru.scala 212:30]
    io_wbreq_wdata2_REG <= s2_out[31:0]; // @[coru.scala 214:36]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_valid <= 1'h0;
    end else if (_T_22) begin
      s1_uop_valid <= io_uopin_valid;
    end else if (flop) begin
      s1_uop_valid <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_cortype <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_cortype <= io_uopin_bits_cortype;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_valid <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_valid <= io_uopin_bits_srcreq_0_valid;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_valid <= s1_uop_bits_srcreq_0_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_idx <= 6'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_idx <= io_uopin_bits_srcreq_0_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_busy <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_busy <= io_uopin_bits_srcreq_0_busy;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_busy <= s1_uop_bits_srcreq_0_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_0 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_wkupidx_0 <= io_uopin_bits_srcreq_0_wkupidx_0;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_wkupidx_0 <= s1_uop_bits_srcreq_0_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_1 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_wkupidx_1 <= io_uopin_bits_srcreq_0_wkupidx_1;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_wkupidx_1 <= s1_uop_bits_srcreq_0_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_2 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_wkupidx_2 <= io_uopin_bits_srcreq_0_wkupidx_2;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_wkupidx_2 <= s1_uop_bits_srcreq_0_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_3 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_wkupidx_3 <= io_uopin_bits_srcreq_0_wkupidx_3;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_wkupidx_3 <= s1_uop_bits_srcreq_0_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_4 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_wkupidx_4 <= io_uopin_bits_srcreq_0_wkupidx_4;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_wkupidx_4 <= s1_uop_bits_srcreq_0_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_0_wkupidx_5 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_0_wkupidx_5 <= io_uopin_bits_srcreq_0_wkupidx_5;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_0_wkupidx_5 <= s1_uop_bits_srcreq_0_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_valid <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_valid <= io_uopin_bits_srcreq_1_valid;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_valid <= s1_uop_bits_srcreq_1_out_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_idx <= 6'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_idx <= io_uopin_bits_srcreq_1_idx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_busy <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_busy <= io_uopin_bits_srcreq_1_busy;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_busy <= s1_uop_bits_srcreq_1_out_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_0 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_wkupidx_0 <= io_uopin_bits_srcreq_1_wkupidx_0;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_wkupidx_0 <= s1_uop_bits_srcreq_1_out_wkupidx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_1 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_wkupidx_1 <= io_uopin_bits_srcreq_1_wkupidx_1;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_wkupidx_1 <= s1_uop_bits_srcreq_1_out_wkupidx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_2 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_wkupidx_2 <= io_uopin_bits_srcreq_1_wkupidx_2;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_wkupidx_2 <= s1_uop_bits_srcreq_1_out_wkupidx_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_3 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_wkupidx_3 <= io_uopin_bits_srcreq_1_wkupidx_3;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_wkupidx_3 <= s1_uop_bits_srcreq_1_out_wkupidx_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_4 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_wkupidx_4 <= io_uopin_bits_srcreq_1_wkupidx_4;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_wkupidx_4 <= s1_uop_bits_srcreq_1_out_wkupidx_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_srcreq_1_wkupidx_5 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_srcreq_1_wkupidx_5 <= io_uopin_bits_srcreq_1_wkupidx_5;
    end else if (s1_uop_valid) begin
      s1_uop_bits_srcreq_1_wkupidx_5 <= s1_uop_bits_srcreq_1_out_wkupidx_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wbvld <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_wbvld <= io_uopin_bits_wbvld;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wbreq <= 6'h0;
    end else if (_T_22) begin
      s1_uop_bits_wbreq <= io_uopin_bits_wbreq;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_0 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_waridx_0 <= io_uopin_bits_waridx_0;
    end else if (s1_uop_valid) begin
      s1_uop_bits_waridx_0 <= out__0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_1 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_waridx_1 <= io_uopin_bits_waridx_1;
    end else if (s1_uop_valid) begin
      s1_uop_bits_waridx_1 <= out__1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_2 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_waridx_2 <= io_uopin_bits_waridx_2;
    end else if (s1_uop_valid) begin
      s1_uop_bits_waridx_2 <= out__2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_3 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_waridx_3 <= io_uopin_bits_waridx_3;
    end else if (s1_uop_valid) begin
      s1_uop_bits_waridx_3 <= out__3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_waridx_4 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_waridx_4 <= io_uopin_bits_waridx_4;
    end else if (s1_uop_valid) begin
      s1_uop_bits_waridx_4 <= out__4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_0 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_wawidx_0 <= io_uopin_bits_wawidx_0;
    end else if (s1_uop_valid) begin
      s1_uop_bits_wawidx_0 <= out_1_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_1 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_wawidx_1 <= io_uopin_bits_wawidx_1;
    end else if (s1_uop_valid) begin
      s1_uop_bits_wawidx_1 <= out_1_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_2 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_wawidx_2 <= io_uopin_bits_wawidx_2;
    end else if (s1_uop_valid) begin
      s1_uop_bits_wawidx_2 <= out_1_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_3 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_wawidx_3 <= io_uopin_bits_wawidx_3;
    end else if (s1_uop_valid) begin
      s1_uop_bits_wawidx_3 <= out_1_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_uop_bits_wawidx_4 <= 1'h0;
    end else if (_T_22) begin
      s1_uop_bits_wawidx_4 <= io_uopin_bits_wawidx_4;
    end else if (s1_uop_valid) begin
      s1_uop_bits_wawidx_4 <= out_1_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_vld <= 1'h0;
    end else begin
      s2_vld <= s1_uop_valid & flop;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_wbidx <= 6'h0;
    end else begin
      s2_wbidx <= s1_uop_bits_wbreq;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s2_cortype <= 1'h0;
    end else if (_s2_vld_T) begin
      s2_cortype <= s1_uop_bits_cortype;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_data_reg_0 <= 37'sh0;
    end else if (_s2_vld_T) begin
      s1_data_reg_0 <= s1_data_5_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_data_reg_1 <= 37'sh0;
    end else if (_s2_vld_T) begin
      s1_data_reg_1 <= s1_data_5_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      s1_data_reg_2 <= 37'sh0;
    end else if (_s2_vld_T) begin
      s1_data_reg_2 <= s1_data_5_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_uop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s1_uop_bits_cortype = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_idx = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_busy = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  s1_uop_bits_srcreq_0_wkupidx_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_idx = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_busy = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_4 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  s1_uop_bits_srcreq_1_wkupidx_5 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  s1_uop_bits_wbvld = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s1_uop_bits_wbreq = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  s1_uop_bits_waridx_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  s1_uop_bits_waridx_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  s1_uop_bits_waridx_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s1_uop_bits_waridx_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  s1_uop_bits_waridx_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  s1_uop_bits_wawidx_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  s1_uop_bits_wawidx_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  s1_uop_bits_wawidx_2 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  s1_uop_bits_wawidx_3 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  s1_uop_bits_wawidx_4 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  s2_vld = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  s2_wbidx = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  s2_cortype = _RAND_34[0:0];
  _RAND_35 = {2{`RANDOM}};
  s1_data_reg_0 = _RAND_35[36:0];
  _RAND_36 = {2{`RANDOM}};
  s1_data_reg_1 = _RAND_36[36:0];
  _RAND_37 = {2{`RANDOM}};
  s1_data_reg_2 = _RAND_37[36:0];
  _RAND_38 = {1{`RANDOM}};
  io_wbreq_vld_REG = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  io_wbreq_gregidx_REG = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  io_wbreq_wdata2_REG = _RAND_40[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    s1_uop_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_cortype = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_0_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_valid = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_idx = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_busy = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_srcreq_1_wkupidx_5 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wbvld = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wbreq = 6'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_waridx_4 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_0 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_1 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_2 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_3 = 1'h0;
  end
  if (reset) begin
    s1_uop_bits_wawidx_4 = 1'h0;
  end
  if (reset) begin
    s2_vld = 1'h0;
  end
  if (reset) begin
    s2_wbidx = 6'h0;
  end
  if (reset) begin
    s2_cortype = 1'h0;
  end
  if (reset) begin
    s1_data_reg_0 = 37'sh0;
  end
  if (reset) begin
    s1_data_reg_1 = 37'sh0;
  end
  if (reset) begin
    s1_data_reg_2 = 37'sh0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DspTop(
  input          clock,
  input          reset,
  output         io_din_ready,
  input          io_din_valid,
  input  [31:0]  io_din_bits_0,
  input  [31:0]  io_din_bits_1,
  input          io_dout_ready,
  output         io_dout_valid,
  output [31:0]  io_dout_bits_0,
  output [31:0]  io_dout_bits_1,
  input          io_coefin_regmap_mainch_alp_en,
  input  [31:0]  io_coefin_regmap_mainch_pre_scale,
  input  [31:0]  io_coefin_regmap_mainch_post_scale,
  input  [287:0] io_coefin_regmap_mainch_drc1_coef,
  input          io_coefin_regmap_mainch_drc1_en,
  input  [2:0]   io_coefin_regmap_mainch_ch1_din_sel,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq0_coef,
  input  [127:0] io_coefin_regmap_mainch_ch1_input_mixer,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq1_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq2_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq3_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq4_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq5_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq6_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq7_coef,
  input  [159:0] io_coefin_regmap_mainch_ch1_bq8_coef,
  input  [31:0]  io_coefin_regmap_mainch_ch1_vol_coef,
  input  [95:0]  io_coefin_regmap_mainch_ch1_out_mixer,
  input  [2:0]   io_coefin_regmap_mainch_ch2_din_sel,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq0_coef,
  input  [127:0] io_coefin_regmap_mainch_ch2_input_mixer,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq1_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq2_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq3_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq4_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq5_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq6_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq7_coef,
  input  [159:0] io_coefin_regmap_mainch_ch2_bq8_coef,
  input  [31:0]  io_coefin_regmap_mainch_ch2_vol_coef,
  input  [95:0]  io_coefin_regmap_mainch_ch2_out_mixer,
  input  [31:0]  io_coefin_regmap_subch_vol_coef,
  input  [1:0]   io_coefin_regmap_subch_vol_sel,
  input  [287:0] io_coefin_regmap_subch_drc2_coef,
  input          io_coefin_regmap_subch_drc2_en,
  input  [95:0]  io_coefin_regmap_subch_ch3_input_mixer,
  input  [159:0] io_coefin_regmap_subch_ch3_bq_coef,
  input  [63:0]  io_coefin_regmap_subch_ch4_input_mixer,
  input          io_coefin_regmap_subch_ch4_input_sel,
  input  [159:0] io_coefin_regmap_subch_ch4_bq0_coef,
  input  [159:0] io_coefin_regmap_subch_ch4_bq1_coef
);
  wire  decode_unit_clock; // @[dsptop.scala 86:27]
  wire  decode_unit_reset; // @[dsptop.scala 86:27]
  wire  decode_unit_io_din_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_din_valid; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_din_bits_0; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_din_bits_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_dout_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_dout_valid; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_dout_bits_0; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_dout_bits_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_valid; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_macuio_0_bits_vlen; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_select; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_drc; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_pow; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_loop; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_drcgain; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_drcnum; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_srcreq_0_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_srcreq_1_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_srcreq_2_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_srcreq_3_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_srcreq_4_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_srcreq_5_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_wbvld; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_0_bits_wbreq; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_waridx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_waridx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_waridx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_waridx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_waridx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_wawidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_wawidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_wawidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_wawidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_0_bits_wawidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_valid; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_macuio_1_bits_vlen; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_select; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_drc; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_pow; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_loop; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_drcgain; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_drcnum; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_srcreq_0_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_srcreq_1_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_srcreq_2_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_srcreq_3_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_srcreq_4_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_srcreq_5_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_wbvld; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_1_bits_wbreq; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_waridx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_waridx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_waridx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_waridx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_waridx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_wawidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_wawidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_wawidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_wawidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_1_bits_wawidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_valid; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_macuio_2_bits_vlen; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_select; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_drc; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_pow; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_loop; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_drcgain; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_drcnum; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_srcreq_0_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_srcreq_1_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_srcreq_2_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_srcreq_3_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_srcreq_4_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_srcreq_5_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_wbvld; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_2_bits_wbreq; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_waridx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_waridx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_waridx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_waridx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_waridx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_wawidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_wawidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_wawidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_wawidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_2_bits_wawidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_valid; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_macuio_3_bits_vlen; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_select; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_drc; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_pow; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_loop; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_drcgain; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_drcnum; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_srcreq_0_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_srcreq_1_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_srcreq_2_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_srcreq_3_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_srcreq_4_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_srcreq_5_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_wbvld; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_3_bits_wbreq; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_waridx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_waridx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_waridx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_waridx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_waridx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_wawidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_wawidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_wawidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_wawidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_3_bits_wawidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_valid; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_macuio_4_bits_vlen; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_select; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_drc; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_pow; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_loop; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_drcgain; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_drcnum; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_srcreq_0_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_srcreq_1_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_srcreq_2_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_srcreq_3_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_srcreq_4_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_isgroup; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_iscoef; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_srcreq_5_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_wbvld; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_macuio_4_bits_wbreq; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_waridx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_waridx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_waridx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_waridx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_waridx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_wawidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_wawidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_wawidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_wawidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_macuio_4_bits_wawidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_wd_check_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_wd_check_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_wd_check_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_wd_check_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_wd_check_2_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_wd_check_2_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_wd_check_3_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_wd_check_3_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_wd_check_4_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_wd_check_4_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_wd_check_5_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_wd_check_5_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_0_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_0_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_0_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_0_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_0_2_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_0_2_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_0_3_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_0_3_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_0_4_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_0_4_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_0_5_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_0_5_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_1_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_1_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_1_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_1_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_1_2_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_1_2_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_1_3_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_1_3_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_1_4_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_1_4_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_1_5_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_1_5_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_2_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_2_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_2_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_2_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_2_2_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_2_2_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_2_3_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_2_3_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_2_4_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_2_4_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_2_5_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_2_5_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_3_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_3_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_3_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_3_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_3_2_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_3_2_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_3_3_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_3_3_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_3_4_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_3_4_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_3_5_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_3_5_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_4_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_4_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_4_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_4_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_4_2_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_4_2_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_4_3_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_4_3_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_4_4_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_4_4_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_mac_r_check_4_5_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_mac_r_check_4_5_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_cor_r_check_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_cor_r_check_0_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_cor_r_check_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_cor_r_check_1_bits; // @[dsptop.scala 86:27]
  wire  decode_unit_io_exuempty_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_exuempty_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_exuempty_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_exuempty_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_exuempty_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_exuempty_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_ready; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_valid; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_cortype; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_coruio_bits_srcreq_0_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_valid; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_coruio_bits_srcreq_1_idx; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_busy; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_wbvld; // @[dsptop.scala 86:27]
  wire [5:0] decode_unit_io_coruio_bits_wbreq; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_waridx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_waridx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_waridx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_waridx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_waridx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_wawidx_0; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_wawidx_1; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_wawidx_2; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_wawidx_3; // @[dsptop.scala 86:27]
  wire  decode_unit_io_coruio_bits_wawidx_4; // @[dsptop.scala 86:27]
  wire  decode_unit_io_writerf_valid; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_writerf_bits_0; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_writerf_bits_1; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_writerf_bits_2; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_writerf_bits_3; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_readrf_0; // @[dsptop.scala 86:27]
  wire [31:0] decode_unit_io_readrf_1; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_coef_in_mainch_ch0_inputsel; // @[dsptop.scala 86:27]
  wire [2:0] decode_unit_io_coef_in_mainch_ch1_inputsel; // @[dsptop.scala 86:27]
  wire  reg_file_clock; // @[dsptop.scala 87:27]
  wire  reg_file_reset; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_0_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_0_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_0_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_0_req_gidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_0_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_1_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_1_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_1_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_1_req_gidx; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_1_req_sel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_1_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_2_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_2_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_2_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_2_req_gidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_2_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_3_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_3_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_3_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_3_req_gidx; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_3_req_sel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_3_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_4_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_4_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_4_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_4_req_gidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_4_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_5_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_5_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_5_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_5_req_gidx; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_5_req_sel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_5_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_6_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_6_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_6_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_6_req_gidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_6_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_7_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_7_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_7_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_7_req_gidx; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_7_req_sel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_7_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_8_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_8_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_8_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_8_req_gidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_8_resp; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_9_req_isgroup; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_9_req_iscoef; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_9_req_idx; // @[dsptop.scala 87:27]
  wire [2:0] reg_file_io_exe_rd_9_req_gidx; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_rd_9_req_sel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_9_resp; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_10_req_idx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_10_resp; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_rd_11_req_idx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_rd_11_resp; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_0_wdata1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_0_wdata2; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_wb_0_vld; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_wb_0_gregidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_1_wdata1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_1_wdata2; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_wb_1_vld; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_wb_1_gregidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_2_wdata1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_2_wdata2; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_wb_2_vld; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_wb_2_gregidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_3_wdata1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_3_wdata2; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_wb_3_vld; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_wb_3_gregidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_4_wdata1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_4_wdata2; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_wb_4_vld; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_wb_4_gregidx; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_exe_wb_5_wdata2; // @[dsptop.scala 87:27]
  wire  reg_file_io_exe_wb_5_vld; // @[dsptop.scala 87:27]
  wire [5:0] reg_file_io_exe_wb_5_gregidx; // @[dsptop.scala 87:27]
  wire  reg_file_io_dec_wb_valid; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_dec_wb_bits_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_dec_wb_bits_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_dec_wb_bits_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_dec_wb_bits_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_dec_rd_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_dec_rd_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2mix_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2mix_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2mix_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2bq_0_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2bq_0_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2bq_0_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2bq_0_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2bq_0_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch2vol; // @[dsptop.scala 87:27]
  wire  reg_file_io_coef_in_subch_ch2volsel; // @[dsptop.scala 87:27]
  wire  reg_file_io_coef_in_subch_ch3sel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3mix_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3mix_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_0_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_0_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_0_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_0_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_0_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_1_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_1_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_1_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_1_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3bq_1_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_ch3vol; // @[dsptop.scala 87:27]
  wire  reg_file_io_coef_in_subch_ch3volsel; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_pow_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_pow_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_smooth_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_smooth_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_smooth_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_smooth_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_subch_drc_ratio; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_0_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_0_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_0_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_0_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_0_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_1_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_1_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_1_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_1_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_1_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_2_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_2_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_2_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_2_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_2_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_3_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_3_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_3_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_3_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_3_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_4_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_4_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_4_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_4_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_4_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_5_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_5_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_5_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_5_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_5_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_6_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_6_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_6_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_6_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_6_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_7_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_7_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_7_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_7_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_7_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_8_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_8_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_8_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_8_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_bqcoef_8_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_inputmix_0_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_inputmix_0_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_inputmix_1_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_inputmix_1_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_vol; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_outputmix_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_outputmix_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_outputmix_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_prescale; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch0_postscale; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_0_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_0_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_0_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_0_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_0_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_1_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_1_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_1_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_1_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_1_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_2_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_2_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_2_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_2_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_2_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_3_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_3_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_3_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_3_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_3_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_4_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_4_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_4_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_4_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_4_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_5_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_5_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_5_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_5_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_5_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_6_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_6_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_6_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_6_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_6_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_7_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_7_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_7_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_7_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_7_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_8_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_8_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_8_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_8_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_bqcoef_8_4; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_inputmix_0_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_inputmix_0_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_inputmix_1_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_inputmix_1_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_vol; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_outputmix_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_outputmix_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_ch1_outputmix_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_pow_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_pow_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_smooth_0; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_smooth_1; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_smooth_2; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_smooth_3; // @[dsptop.scala 87:27]
  wire [31:0] reg_file_io_coef_in_mainch_drc_ratio; // @[dsptop.scala 87:27]
  wire  mac_units_0_clock; // @[dsptop.scala 88:70]
  wire  mac_units_0_reset; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_ready; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_valid; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_0_io_uopin_bits_vlen; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_select; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_drc; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_pow; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_loop; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_drcgain; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_drcnum; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_valid; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_srcreq_0_idx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_busy; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_valid; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_srcreq_1_idx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_busy; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_valid; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_srcreq_2_idx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_busy; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_valid; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_srcreq_3_idx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_busy; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_valid; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_srcreq_4_idx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_busy; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_valid; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_srcreq_5_idx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_busy; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_wbvld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_uopin_bits_wbreq; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_waridx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_waridx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_waridx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_waridx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_waridx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_wawidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_wawidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_wawidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_wawidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_uopin_bits_wawidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_rfreq_0_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_rfreq_0_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_rfreq_0_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_0_io_rfreq_0_req_gidx; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_rfreq_0_resp; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_rfreq_1_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_rfreq_1_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_rfreq_1_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_0_io_rfreq_1_req_gidx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_rfreq_1_req_sel; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_rfreq_1_resp; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_wbreq_wdata1; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_wbreq_wdata2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_wbreq_vld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_wbreq_gregidx; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_empty; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_raw_wkup_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_raw_wkup_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_raw_wkup_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_raw_wkup_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_raw_wkup_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_raw_wkup_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_raw_wkup_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_raw_wkup_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_raw_wkup_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_raw_wkup_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_raw_wkup_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_raw_wkup_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_wbcheck_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_wbcheck_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_r_check_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_r_check_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_r_check_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_r_check_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_r_check_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_r_check_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_r_check_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_r_check_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_r_check_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_r_check_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_r_check_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_0_io_r_check_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_other_flop_0; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_other_flop_1; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_other_flop_2; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_other_flop_3; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_other_flop_4; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_flop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_coef_subch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_coef_subch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_coef_subch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_coef_mainch_ch0_autoloop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_coef_mainch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_0_io_coef_mainch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_0_io_coef_mainch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_1_clock; // @[dsptop.scala 88:70]
  wire  mac_units_1_reset; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_ready; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_valid; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_1_io_uopin_bits_vlen; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_select; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_drc; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_pow; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_loop; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_drcgain; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_drcnum; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_valid; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_srcreq_0_idx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_busy; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_valid; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_srcreq_1_idx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_busy; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_valid; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_srcreq_2_idx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_busy; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_valid; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_srcreq_3_idx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_busy; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_valid; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_srcreq_4_idx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_busy; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_valid; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_srcreq_5_idx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_busy; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_wbvld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_uopin_bits_wbreq; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_waridx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_waridx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_waridx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_waridx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_waridx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_wawidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_wawidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_wawidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_wawidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_uopin_bits_wawidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_rfreq_0_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_rfreq_0_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_rfreq_0_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_1_io_rfreq_0_req_gidx; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_rfreq_0_resp; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_rfreq_1_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_rfreq_1_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_rfreq_1_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_1_io_rfreq_1_req_gidx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_rfreq_1_req_sel; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_rfreq_1_resp; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_wbreq_wdata1; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_wbreq_wdata2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_wbreq_vld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_wbreq_gregidx; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_empty; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_raw_wkup_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_raw_wkup_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_raw_wkup_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_raw_wkup_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_raw_wkup_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_raw_wkup_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_raw_wkup_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_raw_wkup_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_raw_wkup_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_raw_wkup_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_raw_wkup_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_raw_wkup_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_wbcheck_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_wbcheck_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_r_check_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_r_check_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_r_check_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_r_check_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_r_check_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_r_check_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_r_check_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_r_check_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_r_check_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_r_check_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_r_check_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_1_io_r_check_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_other_flop_0; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_other_flop_1; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_other_flop_2; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_other_flop_3; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_other_flop_4; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_flop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_coef_subch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_coef_subch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_coef_subch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_coef_mainch_ch0_autoloop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_coef_mainch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_1_io_coef_mainch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_1_io_coef_mainch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_2_clock; // @[dsptop.scala 88:70]
  wire  mac_units_2_reset; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_ready; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_valid; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_2_io_uopin_bits_vlen; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_select; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_drc; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_pow; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_loop; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_drcgain; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_drcnum; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_valid; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_srcreq_0_idx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_busy; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_valid; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_srcreq_1_idx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_busy; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_valid; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_srcreq_2_idx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_busy; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_valid; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_srcreq_3_idx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_busy; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_valid; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_srcreq_4_idx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_busy; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_valid; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_srcreq_5_idx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_busy; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_wbvld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_uopin_bits_wbreq; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_waridx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_waridx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_waridx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_waridx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_waridx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_wawidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_wawidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_wawidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_wawidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_uopin_bits_wawidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_rfreq_0_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_rfreq_0_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_rfreq_0_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_2_io_rfreq_0_req_gidx; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_rfreq_0_resp; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_rfreq_1_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_rfreq_1_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_rfreq_1_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_2_io_rfreq_1_req_gidx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_rfreq_1_req_sel; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_rfreq_1_resp; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_wbreq_wdata1; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_wbreq_wdata2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_wbreq_vld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_wbreq_gregidx; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_empty; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_raw_wkup_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_raw_wkup_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_raw_wkup_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_raw_wkup_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_raw_wkup_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_raw_wkup_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_raw_wkup_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_raw_wkup_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_raw_wkup_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_raw_wkup_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_raw_wkup_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_raw_wkup_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_wbcheck_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_wbcheck_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_r_check_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_r_check_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_r_check_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_r_check_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_r_check_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_r_check_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_r_check_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_r_check_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_r_check_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_r_check_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_r_check_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_2_io_r_check_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_other_flop_0; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_other_flop_1; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_other_flop_2; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_other_flop_3; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_other_flop_4; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_flop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_coef_subch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_coef_subch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_coef_subch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_coef_mainch_ch0_autoloop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_coef_mainch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_2_io_coef_mainch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_2_io_coef_mainch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_3_clock; // @[dsptop.scala 88:70]
  wire  mac_units_3_reset; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_ready; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_valid; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_3_io_uopin_bits_vlen; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_select; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_drc; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_pow; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_loop; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_drcgain; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_drcnum; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_valid; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_srcreq_0_idx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_busy; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_valid; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_srcreq_1_idx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_busy; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_valid; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_srcreq_2_idx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_busy; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_valid; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_srcreq_3_idx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_busy; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_valid; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_srcreq_4_idx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_busy; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_valid; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_srcreq_5_idx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_busy; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_wbvld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_uopin_bits_wbreq; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_waridx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_waridx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_waridx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_waridx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_waridx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_wawidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_wawidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_wawidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_wawidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_uopin_bits_wawidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_rfreq_0_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_rfreq_0_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_rfreq_0_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_3_io_rfreq_0_req_gidx; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_rfreq_0_resp; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_rfreq_1_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_rfreq_1_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_rfreq_1_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_3_io_rfreq_1_req_gidx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_rfreq_1_req_sel; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_rfreq_1_resp; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_wbreq_wdata1; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_wbreq_wdata2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_wbreq_vld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_wbreq_gregidx; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_empty; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_raw_wkup_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_raw_wkup_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_raw_wkup_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_raw_wkup_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_raw_wkup_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_raw_wkup_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_raw_wkup_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_raw_wkup_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_raw_wkup_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_raw_wkup_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_raw_wkup_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_raw_wkup_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_wbcheck_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_wbcheck_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_r_check_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_r_check_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_r_check_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_r_check_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_r_check_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_r_check_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_r_check_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_r_check_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_r_check_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_r_check_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_r_check_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_3_io_r_check_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_other_flop_0; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_other_flop_1; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_other_flop_2; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_other_flop_3; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_other_flop_4; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_flop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_coef_subch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_coef_subch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_coef_subch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_coef_mainch_ch0_autoloop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_coef_mainch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_3_io_coef_mainch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_3_io_coef_mainch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_4_clock; // @[dsptop.scala 88:70]
  wire  mac_units_4_reset; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_ready; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_valid; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_4_io_uopin_bits_vlen; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_select; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_drc; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_pow; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_loop; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_drcgain; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_drcnum; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_valid; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_srcreq_0_idx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_busy; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_valid; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_srcreq_1_idx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_busy; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_valid; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_srcreq_2_idx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_busy; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_valid; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_srcreq_3_idx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_busy; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_valid; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_srcreq_4_idx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_busy; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_valid; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_srcreq_5_idx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_busy; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_wbvld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_uopin_bits_wbreq; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_waridx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_waridx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_waridx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_waridx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_waridx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_wawidx_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_wawidx_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_wawidx_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_wawidx_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_uopin_bits_wawidx_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_rfreq_0_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_rfreq_0_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_rfreq_0_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_4_io_rfreq_0_req_gidx; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_rfreq_0_resp; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_rfreq_1_req_isgroup; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_rfreq_1_req_iscoef; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_rfreq_1_req_idx; // @[dsptop.scala 88:70]
  wire [2:0] mac_units_4_io_rfreq_1_req_gidx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_rfreq_1_req_sel; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_rfreq_1_resp; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_wbreq_wdata1; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_wbreq_wdata2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_wbreq_vld; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_wbreq_gregidx; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_empty; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_raw_wkup_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_raw_wkup_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_raw_wkup_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_raw_wkup_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_raw_wkup_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_raw_wkup_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_raw_wkup_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_raw_wkup_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_raw_wkup_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_raw_wkup_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_raw_wkup_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_raw_wkup_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_wbcheck_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_wbcheck_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_r_check_0_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_r_check_0_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_r_check_1_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_r_check_1_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_r_check_2_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_r_check_2_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_r_check_3_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_r_check_3_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_r_check_4_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_r_check_4_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_r_check_5_valid; // @[dsptop.scala 88:70]
  wire [5:0] mac_units_4_io_r_check_5_bits; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_other_flop_0; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_other_flop_1; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_other_flop_2; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_other_flop_3; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_other_flop_4; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_flop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_coef_subch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_coef_subch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_coef_subch_drc_drcen; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_coef_mainch_ch0_autoloop; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_coef_mainch_drc_th; // @[dsptop.scala 88:70]
  wire [31:0] mac_units_4_io_coef_mainch_drc_offset; // @[dsptop.scala 88:70]
  wire  mac_units_4_io_coef_mainch_drc_drcen; // @[dsptop.scala 88:70]
  wire  cor_unit_clock; // @[dsptop.scala 89:27]
  wire  cor_unit_reset; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_ready; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_valid; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_cortype; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_uopin_bits_srcreq_0_idx; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_busy; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_uopin_bits_srcreq_1_idx; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_busy; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_wbvld; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_uopin_bits_wbreq; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_waridx_0; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_waridx_1; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_waridx_2; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_waridx_3; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_waridx_4; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_wawidx_0; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_wawidx_1; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_wawidx_2; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_wawidx_3; // @[dsptop.scala 89:27]
  wire  cor_unit_io_uopin_bits_wawidx_4; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_rfreq_0_req_idx; // @[dsptop.scala 89:27]
  wire [31:0] cor_unit_io_rfreq_0_resp; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_rfreq_1_req_idx; // @[dsptop.scala 89:27]
  wire [31:0] cor_unit_io_rfreq_1_resp; // @[dsptop.scala 89:27]
  wire [31:0] cor_unit_io_wbreq_wdata2; // @[dsptop.scala 89:27]
  wire  cor_unit_io_wbreq_vld; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_wbreq_gregidx; // @[dsptop.scala 89:27]
  wire  cor_unit_io_empty; // @[dsptop.scala 89:27]
  wire  cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_raw_wkup_0_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_raw_wkup_0_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_raw_wkup_1_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_raw_wkup_1_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_raw_wkup_2_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_raw_wkup_2_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_raw_wkup_3_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_raw_wkup_3_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_raw_wkup_4_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_raw_wkup_4_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_raw_wkup_5_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_raw_wkup_5_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_wbcheck_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_wbcheck_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_r_check_0_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_r_check_0_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_r_check_1_valid; // @[dsptop.scala 89:27]
  wire [5:0] cor_unit_io_r_check_1_bits; // @[dsptop.scala 89:27]
  wire  cor_unit_io_other_flop_0; // @[dsptop.scala 89:27]
  wire  cor_unit_io_other_flop_1; // @[dsptop.scala 89:27]
  wire  cor_unit_io_other_flop_2; // @[dsptop.scala 89:27]
  wire  cor_unit_io_other_flop_3; // @[dsptop.scala 89:27]
  wire  cor_unit_io_other_flop_4; // @[dsptop.scala 89:27]
  wire  cor_unit_io_flop; // @[dsptop.scala 89:27]
  wire [5:0] coef_mainch_drc_pow_0_hi = io_coefin_regmap_mainch_drc1_coef[281] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_pow_0_lo = io_coefin_regmap_mainch_drc1_coef[281:256]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_pow_1_hi = io_coefin_regmap_mainch_drc1_coef[249] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_pow_1_lo = io_coefin_regmap_mainch_drc1_coef[249:224]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_smooth_0_hi = io_coefin_regmap_mainch_drc1_coef[217] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_smooth_0_lo = io_coefin_regmap_mainch_drc1_coef[217:192]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_smooth_1_hi = io_coefin_regmap_mainch_drc1_coef[185] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_smooth_1_lo = io_coefin_regmap_mainch_drc1_coef[185:160]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_smooth_2_hi = io_coefin_regmap_mainch_drc1_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_smooth_2_lo = io_coefin_regmap_mainch_drc1_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_smooth_3_hi = io_coefin_regmap_mainch_drc1_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_smooth_3_lo = io_coefin_regmap_mainch_drc1_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_ratio_hi = io_coefin_regmap_mainch_drc1_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_ratio_lo = io_coefin_regmap_mainch_drc1_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_drc_offset_hi = io_coefin_regmap_mainch_drc1_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_drc_offset_lo = io_coefin_regmap_mainch_drc1_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_pow_0_hi = io_coefin_regmap_subch_drc2_coef[281] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_pow_0_lo = io_coefin_regmap_subch_drc2_coef[281:256]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_pow_1_hi = io_coefin_regmap_subch_drc2_coef[249] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_pow_1_lo = io_coefin_regmap_subch_drc2_coef[249:224]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_smooth_0_hi = io_coefin_regmap_subch_drc2_coef[217] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_smooth_0_lo = io_coefin_regmap_subch_drc2_coef[217:192]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_smooth_1_hi = io_coefin_regmap_subch_drc2_coef[185] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_smooth_1_lo = io_coefin_regmap_subch_drc2_coef[185:160]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_smooth_2_hi = io_coefin_regmap_subch_drc2_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_smooth_2_lo = io_coefin_regmap_subch_drc2_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_smooth_3_hi = io_coefin_regmap_subch_drc2_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_smooth_3_lo = io_coefin_regmap_subch_drc2_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_ratio_hi = io_coefin_regmap_subch_drc2_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_ratio_lo = io_coefin_regmap_subch_drc2_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_drc_offset_hi = io_coefin_regmap_subch_drc2_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_drc_offset_lo = io_coefin_regmap_subch_drc2_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_postscale_hi = io_coefin_regmap_mainch_post_scale[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_postscale_lo = io_coefin_regmap_mainch_post_scale[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_0_0_hi = io_coefin_regmap_mainch_ch1_bq0_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_0_0_lo = io_coefin_regmap_mainch_ch1_bq0_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_0_1_hi = io_coefin_regmap_mainch_ch1_bq0_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_0_1_lo = io_coefin_regmap_mainch_ch1_bq0_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_0_2_hi = io_coefin_regmap_mainch_ch1_bq0_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_0_2_lo = io_coefin_regmap_mainch_ch1_bq0_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_0_3_hi = io_coefin_regmap_mainch_ch1_bq0_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_0_3_lo = io_coefin_regmap_mainch_ch1_bq0_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_0_4_hi = io_coefin_regmap_mainch_ch1_bq0_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_0_4_lo = io_coefin_regmap_mainch_ch1_bq0_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_1_0_hi = io_coefin_regmap_mainch_ch1_bq1_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_1_0_lo = io_coefin_regmap_mainch_ch1_bq1_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_1_1_hi = io_coefin_regmap_mainch_ch1_bq1_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_1_1_lo = io_coefin_regmap_mainch_ch1_bq1_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_1_2_hi = io_coefin_regmap_mainch_ch1_bq1_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_1_2_lo = io_coefin_regmap_mainch_ch1_bq1_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_1_3_hi = io_coefin_regmap_mainch_ch1_bq1_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_1_3_lo = io_coefin_regmap_mainch_ch1_bq1_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_1_4_hi = io_coefin_regmap_mainch_ch1_bq1_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_1_4_lo = io_coefin_regmap_mainch_ch1_bq1_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_2_0_hi = io_coefin_regmap_mainch_ch1_bq2_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_2_0_lo = io_coefin_regmap_mainch_ch1_bq2_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_2_1_hi = io_coefin_regmap_mainch_ch1_bq2_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_2_1_lo = io_coefin_regmap_mainch_ch1_bq2_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_2_2_hi = io_coefin_regmap_mainch_ch1_bq2_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_2_2_lo = io_coefin_regmap_mainch_ch1_bq2_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_2_3_hi = io_coefin_regmap_mainch_ch1_bq2_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_2_3_lo = io_coefin_regmap_mainch_ch1_bq2_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_2_4_hi = io_coefin_regmap_mainch_ch1_bq2_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_2_4_lo = io_coefin_regmap_mainch_ch1_bq2_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_3_0_hi = io_coefin_regmap_mainch_ch1_bq3_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_3_0_lo = io_coefin_regmap_mainch_ch1_bq3_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_3_1_hi = io_coefin_regmap_mainch_ch1_bq3_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_3_1_lo = io_coefin_regmap_mainch_ch1_bq3_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_3_2_hi = io_coefin_regmap_mainch_ch1_bq3_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_3_2_lo = io_coefin_regmap_mainch_ch1_bq3_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_3_3_hi = io_coefin_regmap_mainch_ch1_bq3_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_3_3_lo = io_coefin_regmap_mainch_ch1_bq3_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_3_4_hi = io_coefin_regmap_mainch_ch1_bq3_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_3_4_lo = io_coefin_regmap_mainch_ch1_bq3_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_4_0_hi = io_coefin_regmap_mainch_ch1_bq4_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_4_0_lo = io_coefin_regmap_mainch_ch1_bq4_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_4_1_hi = io_coefin_regmap_mainch_ch1_bq4_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_4_1_lo = io_coefin_regmap_mainch_ch1_bq4_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_4_2_hi = io_coefin_regmap_mainch_ch1_bq4_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_4_2_lo = io_coefin_regmap_mainch_ch1_bq4_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_4_3_hi = io_coefin_regmap_mainch_ch1_bq4_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_4_3_lo = io_coefin_regmap_mainch_ch1_bq4_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_4_4_hi = io_coefin_regmap_mainch_ch1_bq4_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_4_4_lo = io_coefin_regmap_mainch_ch1_bq4_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_5_0_hi = io_coefin_regmap_mainch_ch1_bq5_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_5_0_lo = io_coefin_regmap_mainch_ch1_bq5_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_5_1_hi = io_coefin_regmap_mainch_ch1_bq5_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_5_1_lo = io_coefin_regmap_mainch_ch1_bq5_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_5_2_hi = io_coefin_regmap_mainch_ch1_bq5_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_5_2_lo = io_coefin_regmap_mainch_ch1_bq5_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_5_3_hi = io_coefin_regmap_mainch_ch1_bq5_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_5_3_lo = io_coefin_regmap_mainch_ch1_bq5_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_5_4_hi = io_coefin_regmap_mainch_ch1_bq5_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_5_4_lo = io_coefin_regmap_mainch_ch1_bq5_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_6_0_hi = io_coefin_regmap_mainch_ch1_bq6_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_6_0_lo = io_coefin_regmap_mainch_ch1_bq6_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_6_1_hi = io_coefin_regmap_mainch_ch1_bq6_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_6_1_lo = io_coefin_regmap_mainch_ch1_bq6_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_6_2_hi = io_coefin_regmap_mainch_ch1_bq6_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_6_2_lo = io_coefin_regmap_mainch_ch1_bq6_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_6_3_hi = io_coefin_regmap_mainch_ch1_bq6_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_6_3_lo = io_coefin_regmap_mainch_ch1_bq6_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_6_4_hi = io_coefin_regmap_mainch_ch1_bq6_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_6_4_lo = io_coefin_regmap_mainch_ch1_bq6_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_7_0_hi = io_coefin_regmap_mainch_ch1_bq7_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_7_0_lo = io_coefin_regmap_mainch_ch1_bq7_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_7_1_hi = io_coefin_regmap_mainch_ch1_bq7_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_7_1_lo = io_coefin_regmap_mainch_ch1_bq7_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_7_2_hi = io_coefin_regmap_mainch_ch1_bq7_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_7_2_lo = io_coefin_regmap_mainch_ch1_bq7_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_7_3_hi = io_coefin_regmap_mainch_ch1_bq7_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_7_3_lo = io_coefin_regmap_mainch_ch1_bq7_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_7_4_hi = io_coefin_regmap_mainch_ch1_bq7_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_7_4_lo = io_coefin_regmap_mainch_ch1_bq7_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_8_0_hi = io_coefin_regmap_mainch_ch1_bq8_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_8_0_lo = io_coefin_regmap_mainch_ch1_bq8_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_8_1_hi = io_coefin_regmap_mainch_ch1_bq8_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_8_1_lo = io_coefin_regmap_mainch_ch1_bq8_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_8_2_hi = io_coefin_regmap_mainch_ch1_bq8_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_8_2_lo = io_coefin_regmap_mainch_ch1_bq8_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_8_3_hi = io_coefin_regmap_mainch_ch1_bq8_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_8_3_lo = io_coefin_regmap_mainch_ch1_bq8_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_bqcoef_8_4_hi = io_coefin_regmap_mainch_ch1_bq8_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_bqcoef_8_4_lo = io_coefin_regmap_mainch_ch1_bq8_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_outputmix_0_hi = io_coefin_regmap_mainch_ch1_out_mixer[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_outputmix_0_lo = io_coefin_regmap_mainch_ch1_out_mixer[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_outputmix_1_hi = io_coefin_regmap_mainch_ch1_out_mixer[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_outputmix_1_lo = io_coefin_regmap_mainch_ch1_out_mixer[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_outputmix_2_hi = io_coefin_regmap_mainch_ch1_out_mixer[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_outputmix_2_lo = io_coefin_regmap_mainch_ch1_out_mixer[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_inputmix_0_0_hi = io_coefin_regmap_mainch_ch1_input_mixer[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_inputmix_0_0_lo = io_coefin_regmap_mainch_ch1_input_mixer[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_inputmix_0_1_hi = io_coefin_regmap_mainch_ch1_input_mixer[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_inputmix_0_1_lo = io_coefin_regmap_mainch_ch1_input_mixer[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_inputmix_1_0_hi = io_coefin_regmap_mainch_ch1_input_mixer[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_inputmix_1_0_lo = io_coefin_regmap_mainch_ch1_input_mixer[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch0_inputmix_1_1_hi = io_coefin_regmap_mainch_ch1_input_mixer[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch0_inputmix_1_1_lo = io_coefin_regmap_mainch_ch1_input_mixer[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_0_0_hi = io_coefin_regmap_mainch_ch2_bq0_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_0_0_lo = io_coefin_regmap_mainch_ch2_bq0_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_0_1_hi = io_coefin_regmap_mainch_ch2_bq0_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_0_1_lo = io_coefin_regmap_mainch_ch2_bq0_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_0_2_hi = io_coefin_regmap_mainch_ch2_bq0_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_0_2_lo = io_coefin_regmap_mainch_ch2_bq0_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_0_3_hi = io_coefin_regmap_mainch_ch2_bq0_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_0_3_lo = io_coefin_regmap_mainch_ch2_bq0_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_0_4_hi = io_coefin_regmap_mainch_ch2_bq0_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_0_4_lo = io_coefin_regmap_mainch_ch2_bq0_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_1_0_hi = io_coefin_regmap_mainch_ch2_bq1_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_1_0_lo = io_coefin_regmap_mainch_ch2_bq1_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_1_1_hi = io_coefin_regmap_mainch_ch2_bq1_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_1_1_lo = io_coefin_regmap_mainch_ch2_bq1_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_1_2_hi = io_coefin_regmap_mainch_ch2_bq1_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_1_2_lo = io_coefin_regmap_mainch_ch2_bq1_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_1_3_hi = io_coefin_regmap_mainch_ch2_bq1_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_1_3_lo = io_coefin_regmap_mainch_ch2_bq1_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_1_4_hi = io_coefin_regmap_mainch_ch2_bq1_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_1_4_lo = io_coefin_regmap_mainch_ch2_bq1_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_2_0_hi = io_coefin_regmap_mainch_ch2_bq2_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_2_0_lo = io_coefin_regmap_mainch_ch2_bq2_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_2_1_hi = io_coefin_regmap_mainch_ch2_bq2_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_2_1_lo = io_coefin_regmap_mainch_ch2_bq2_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_2_2_hi = io_coefin_regmap_mainch_ch2_bq2_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_2_2_lo = io_coefin_regmap_mainch_ch2_bq2_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_2_3_hi = io_coefin_regmap_mainch_ch2_bq2_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_2_3_lo = io_coefin_regmap_mainch_ch2_bq2_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_2_4_hi = io_coefin_regmap_mainch_ch2_bq2_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_2_4_lo = io_coefin_regmap_mainch_ch2_bq2_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_3_0_hi = io_coefin_regmap_mainch_ch2_bq3_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_3_0_lo = io_coefin_regmap_mainch_ch2_bq3_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_3_1_hi = io_coefin_regmap_mainch_ch2_bq3_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_3_1_lo = io_coefin_regmap_mainch_ch2_bq3_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_3_2_hi = io_coefin_regmap_mainch_ch2_bq3_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_3_2_lo = io_coefin_regmap_mainch_ch2_bq3_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_3_3_hi = io_coefin_regmap_mainch_ch2_bq3_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_3_3_lo = io_coefin_regmap_mainch_ch2_bq3_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_3_4_hi = io_coefin_regmap_mainch_ch2_bq3_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_3_4_lo = io_coefin_regmap_mainch_ch2_bq3_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_4_0_hi = io_coefin_regmap_mainch_ch2_bq4_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_4_0_lo = io_coefin_regmap_mainch_ch2_bq4_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_4_1_hi = io_coefin_regmap_mainch_ch2_bq4_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_4_1_lo = io_coefin_regmap_mainch_ch2_bq4_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_4_2_hi = io_coefin_regmap_mainch_ch2_bq4_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_4_2_lo = io_coefin_regmap_mainch_ch2_bq4_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_4_3_hi = io_coefin_regmap_mainch_ch2_bq4_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_4_3_lo = io_coefin_regmap_mainch_ch2_bq4_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_4_4_hi = io_coefin_regmap_mainch_ch2_bq4_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_4_4_lo = io_coefin_regmap_mainch_ch2_bq4_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_5_0_hi = io_coefin_regmap_mainch_ch2_bq5_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_5_0_lo = io_coefin_regmap_mainch_ch2_bq5_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_5_1_hi = io_coefin_regmap_mainch_ch2_bq5_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_5_1_lo = io_coefin_regmap_mainch_ch2_bq5_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_5_2_hi = io_coefin_regmap_mainch_ch2_bq5_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_5_2_lo = io_coefin_regmap_mainch_ch2_bq5_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_5_3_hi = io_coefin_regmap_mainch_ch2_bq5_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_5_3_lo = io_coefin_regmap_mainch_ch2_bq5_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_5_4_hi = io_coefin_regmap_mainch_ch2_bq5_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_5_4_lo = io_coefin_regmap_mainch_ch2_bq5_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_6_0_hi = io_coefin_regmap_mainch_ch2_bq6_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_6_0_lo = io_coefin_regmap_mainch_ch2_bq6_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_6_1_hi = io_coefin_regmap_mainch_ch2_bq6_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_6_1_lo = io_coefin_regmap_mainch_ch2_bq6_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_6_2_hi = io_coefin_regmap_mainch_ch2_bq6_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_6_2_lo = io_coefin_regmap_mainch_ch2_bq6_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_6_3_hi = io_coefin_regmap_mainch_ch2_bq6_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_6_3_lo = io_coefin_regmap_mainch_ch2_bq6_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_6_4_hi = io_coefin_regmap_mainch_ch2_bq6_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_6_4_lo = io_coefin_regmap_mainch_ch2_bq6_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_7_0_hi = io_coefin_regmap_mainch_ch2_bq7_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_7_0_lo = io_coefin_regmap_mainch_ch2_bq7_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_7_1_hi = io_coefin_regmap_mainch_ch2_bq7_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_7_1_lo = io_coefin_regmap_mainch_ch2_bq7_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_7_2_hi = io_coefin_regmap_mainch_ch2_bq7_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_7_2_lo = io_coefin_regmap_mainch_ch2_bq7_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_7_3_hi = io_coefin_regmap_mainch_ch2_bq7_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_7_3_lo = io_coefin_regmap_mainch_ch2_bq7_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_7_4_hi = io_coefin_regmap_mainch_ch2_bq7_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_7_4_lo = io_coefin_regmap_mainch_ch2_bq7_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_8_0_hi = io_coefin_regmap_mainch_ch2_bq8_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_8_0_lo = io_coefin_regmap_mainch_ch2_bq8_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_8_1_hi = io_coefin_regmap_mainch_ch2_bq8_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_8_1_lo = io_coefin_regmap_mainch_ch2_bq8_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_8_2_hi = io_coefin_regmap_mainch_ch2_bq8_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_8_2_lo = io_coefin_regmap_mainch_ch2_bq8_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_8_3_hi = io_coefin_regmap_mainch_ch2_bq8_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_8_3_lo = io_coefin_regmap_mainch_ch2_bq8_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_bqcoef_8_4_hi = io_coefin_regmap_mainch_ch2_bq8_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_bqcoef_8_4_lo = io_coefin_regmap_mainch_ch2_bq8_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_outputmix_0_hi = io_coefin_regmap_mainch_ch2_out_mixer[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_outputmix_0_lo = io_coefin_regmap_mainch_ch2_out_mixer[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_outputmix_1_hi = io_coefin_regmap_mainch_ch2_out_mixer[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_outputmix_1_lo = io_coefin_regmap_mainch_ch2_out_mixer[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_outputmix_2_hi = io_coefin_regmap_mainch_ch2_out_mixer[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_outputmix_2_lo = io_coefin_regmap_mainch_ch2_out_mixer[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_inputmix_0_0_hi = io_coefin_regmap_mainch_ch2_input_mixer[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_inputmix_0_0_lo = io_coefin_regmap_mainch_ch2_input_mixer[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_inputmix_0_1_hi = io_coefin_regmap_mainch_ch2_input_mixer[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_inputmix_0_1_lo = io_coefin_regmap_mainch_ch2_input_mixer[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_inputmix_1_0_hi = io_coefin_regmap_mainch_ch2_input_mixer[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_inputmix_1_0_lo = io_coefin_regmap_mainch_ch2_input_mixer[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_mainch_ch1_inputmix_1_1_hi = io_coefin_regmap_mainch_ch2_input_mixer[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_mainch_ch1_inputmix_1_1_lo = io_coefin_regmap_mainch_ch2_input_mixer[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2bq_0_0_hi = io_coefin_regmap_subch_ch3_bq_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2bq_0_0_lo = io_coefin_regmap_subch_ch3_bq_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2bq_0_1_hi = io_coefin_regmap_subch_ch3_bq_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2bq_0_1_lo = io_coefin_regmap_subch_ch3_bq_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2bq_0_2_hi = io_coefin_regmap_subch_ch3_bq_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2bq_0_2_lo = io_coefin_regmap_subch_ch3_bq_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2bq_0_3_hi = io_coefin_regmap_subch_ch3_bq_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2bq_0_3_lo = io_coefin_regmap_subch_ch3_bq_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2bq_0_4_hi = io_coefin_regmap_subch_ch3_bq_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2bq_0_4_lo = io_coefin_regmap_subch_ch3_bq_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2mix_0_hi = io_coefin_regmap_subch_ch3_input_mixer[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2mix_0_lo = io_coefin_regmap_subch_ch3_input_mixer[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2mix_1_hi = io_coefin_regmap_subch_ch3_input_mixer[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2mix_1_lo = io_coefin_regmap_subch_ch3_input_mixer[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch2mix_2_hi = io_coefin_regmap_subch_ch3_input_mixer[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch2mix_2_lo = io_coefin_regmap_subch_ch3_input_mixer[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_0_0_hi = io_coefin_regmap_subch_ch4_bq0_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_0_0_lo = io_coefin_regmap_subch_ch4_bq0_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_0_1_hi = io_coefin_regmap_subch_ch4_bq0_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_0_1_lo = io_coefin_regmap_subch_ch4_bq0_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_0_2_hi = io_coefin_regmap_subch_ch4_bq0_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_0_2_lo = io_coefin_regmap_subch_ch4_bq0_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_0_3_hi = io_coefin_regmap_subch_ch4_bq0_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_0_3_lo = io_coefin_regmap_subch_ch4_bq0_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_0_4_hi = io_coefin_regmap_subch_ch4_bq0_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_0_4_lo = io_coefin_regmap_subch_ch4_bq0_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_1_0_hi = io_coefin_regmap_subch_ch4_bq1_coef[153] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_1_0_lo = io_coefin_regmap_subch_ch4_bq1_coef[153:128]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_1_1_hi = io_coefin_regmap_subch_ch4_bq1_coef[121] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_1_1_lo = io_coefin_regmap_subch_ch4_bq1_coef[121:96]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_1_2_hi = io_coefin_regmap_subch_ch4_bq1_coef[89] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_1_2_lo = io_coefin_regmap_subch_ch4_bq1_coef[89:64]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_1_3_hi = io_coefin_regmap_subch_ch4_bq1_coef[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_1_3_lo = io_coefin_regmap_subch_ch4_bq1_coef[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3bq_1_4_hi = io_coefin_regmap_subch_ch4_bq1_coef[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3bq_1_4_lo = io_coefin_regmap_subch_ch4_bq1_coef[25:0]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3mix_0_hi = io_coefin_regmap_subch_ch4_input_mixer[57] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3mix_0_lo = io_coefin_regmap_subch_ch4_input_mixer[57:32]; // @[dsptop.scala 76:41]
  wire [5:0] coef_subch_ch3mix_1_hi = io_coefin_regmap_subch_ch4_input_mixer[25] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [25:0] coef_subch_ch3mix_1_lo = io_coefin_regmap_subch_ch4_input_mixer[25:0]; // @[dsptop.scala 76:41]
  DspDecode decode_unit ( // @[dsptop.scala 86:27]
    .clock(decode_unit_clock),
    .reset(decode_unit_reset),
    .io_din_ready(decode_unit_io_din_ready),
    .io_din_valid(decode_unit_io_din_valid),
    .io_din_bits_0(decode_unit_io_din_bits_0),
    .io_din_bits_1(decode_unit_io_din_bits_1),
    .io_dout_ready(decode_unit_io_dout_ready),
    .io_dout_valid(decode_unit_io_dout_valid),
    .io_dout_bits_0(decode_unit_io_dout_bits_0),
    .io_dout_bits_1(decode_unit_io_dout_bits_1),
    .io_macuio_0_ready(decode_unit_io_macuio_0_ready),
    .io_macuio_0_valid(decode_unit_io_macuio_0_valid),
    .io_macuio_0_bits_vlen(decode_unit_io_macuio_0_bits_vlen),
    .io_macuio_0_bits_select(decode_unit_io_macuio_0_bits_select),
    .io_macuio_0_bits_drc(decode_unit_io_macuio_0_bits_drc),
    .io_macuio_0_bits_pow(decode_unit_io_macuio_0_bits_pow),
    .io_macuio_0_bits_loop(decode_unit_io_macuio_0_bits_loop),
    .io_macuio_0_bits_drcgain(decode_unit_io_macuio_0_bits_drcgain),
    .io_macuio_0_bits_drcnum(decode_unit_io_macuio_0_bits_drcnum),
    .io_macuio_0_bits_srcreq_0_valid(decode_unit_io_macuio_0_bits_srcreq_0_valid),
    .io_macuio_0_bits_srcreq_0_isgroup(decode_unit_io_macuio_0_bits_srcreq_0_isgroup),
    .io_macuio_0_bits_srcreq_0_iscoef(decode_unit_io_macuio_0_bits_srcreq_0_iscoef),
    .io_macuio_0_bits_srcreq_0_idx(decode_unit_io_macuio_0_bits_srcreq_0_idx),
    .io_macuio_0_bits_srcreq_0_busy(decode_unit_io_macuio_0_bits_srcreq_0_busy),
    .io_macuio_0_bits_srcreq_0_wkupidx_0(decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_0),
    .io_macuio_0_bits_srcreq_0_wkupidx_1(decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_1),
    .io_macuio_0_bits_srcreq_0_wkupidx_2(decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_2),
    .io_macuio_0_bits_srcreq_0_wkupidx_3(decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_3),
    .io_macuio_0_bits_srcreq_0_wkupidx_4(decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_4),
    .io_macuio_0_bits_srcreq_0_wkupidx_5(decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_5),
    .io_macuio_0_bits_srcreq_1_valid(decode_unit_io_macuio_0_bits_srcreq_1_valid),
    .io_macuio_0_bits_srcreq_1_isgroup(decode_unit_io_macuio_0_bits_srcreq_1_isgroup),
    .io_macuio_0_bits_srcreq_1_iscoef(decode_unit_io_macuio_0_bits_srcreq_1_iscoef),
    .io_macuio_0_bits_srcreq_1_idx(decode_unit_io_macuio_0_bits_srcreq_1_idx),
    .io_macuio_0_bits_srcreq_1_busy(decode_unit_io_macuio_0_bits_srcreq_1_busy),
    .io_macuio_0_bits_srcreq_1_wkupidx_0(decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_0),
    .io_macuio_0_bits_srcreq_1_wkupidx_1(decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_1),
    .io_macuio_0_bits_srcreq_1_wkupidx_2(decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_2),
    .io_macuio_0_bits_srcreq_1_wkupidx_3(decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_3),
    .io_macuio_0_bits_srcreq_1_wkupidx_4(decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_4),
    .io_macuio_0_bits_srcreq_1_wkupidx_5(decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_5),
    .io_macuio_0_bits_srcreq_2_valid(decode_unit_io_macuio_0_bits_srcreq_2_valid),
    .io_macuio_0_bits_srcreq_2_isgroup(decode_unit_io_macuio_0_bits_srcreq_2_isgroup),
    .io_macuio_0_bits_srcreq_2_iscoef(decode_unit_io_macuio_0_bits_srcreq_2_iscoef),
    .io_macuio_0_bits_srcreq_2_idx(decode_unit_io_macuio_0_bits_srcreq_2_idx),
    .io_macuio_0_bits_srcreq_2_busy(decode_unit_io_macuio_0_bits_srcreq_2_busy),
    .io_macuio_0_bits_srcreq_2_wkupidx_0(decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_0),
    .io_macuio_0_bits_srcreq_2_wkupidx_1(decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_1),
    .io_macuio_0_bits_srcreq_2_wkupidx_2(decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_2),
    .io_macuio_0_bits_srcreq_2_wkupidx_3(decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_3),
    .io_macuio_0_bits_srcreq_2_wkupidx_4(decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_4),
    .io_macuio_0_bits_srcreq_2_wkupidx_5(decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_5),
    .io_macuio_0_bits_srcreq_3_valid(decode_unit_io_macuio_0_bits_srcreq_3_valid),
    .io_macuio_0_bits_srcreq_3_isgroup(decode_unit_io_macuio_0_bits_srcreq_3_isgroup),
    .io_macuio_0_bits_srcreq_3_iscoef(decode_unit_io_macuio_0_bits_srcreq_3_iscoef),
    .io_macuio_0_bits_srcreq_3_idx(decode_unit_io_macuio_0_bits_srcreq_3_idx),
    .io_macuio_0_bits_srcreq_3_busy(decode_unit_io_macuio_0_bits_srcreq_3_busy),
    .io_macuio_0_bits_srcreq_3_wkupidx_0(decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_0),
    .io_macuio_0_bits_srcreq_3_wkupidx_1(decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_1),
    .io_macuio_0_bits_srcreq_3_wkupidx_2(decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_2),
    .io_macuio_0_bits_srcreq_3_wkupidx_3(decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_3),
    .io_macuio_0_bits_srcreq_3_wkupidx_4(decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_4),
    .io_macuio_0_bits_srcreq_3_wkupidx_5(decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_5),
    .io_macuio_0_bits_srcreq_4_valid(decode_unit_io_macuio_0_bits_srcreq_4_valid),
    .io_macuio_0_bits_srcreq_4_isgroup(decode_unit_io_macuio_0_bits_srcreq_4_isgroup),
    .io_macuio_0_bits_srcreq_4_iscoef(decode_unit_io_macuio_0_bits_srcreq_4_iscoef),
    .io_macuio_0_bits_srcreq_4_idx(decode_unit_io_macuio_0_bits_srcreq_4_idx),
    .io_macuio_0_bits_srcreq_4_busy(decode_unit_io_macuio_0_bits_srcreq_4_busy),
    .io_macuio_0_bits_srcreq_4_wkupidx_0(decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_0),
    .io_macuio_0_bits_srcreq_4_wkupidx_1(decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_1),
    .io_macuio_0_bits_srcreq_4_wkupidx_2(decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_2),
    .io_macuio_0_bits_srcreq_4_wkupidx_3(decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_3),
    .io_macuio_0_bits_srcreq_4_wkupidx_4(decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_4),
    .io_macuio_0_bits_srcreq_4_wkupidx_5(decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_5),
    .io_macuio_0_bits_srcreq_5_valid(decode_unit_io_macuio_0_bits_srcreq_5_valid),
    .io_macuio_0_bits_srcreq_5_isgroup(decode_unit_io_macuio_0_bits_srcreq_5_isgroup),
    .io_macuio_0_bits_srcreq_5_iscoef(decode_unit_io_macuio_0_bits_srcreq_5_iscoef),
    .io_macuio_0_bits_srcreq_5_idx(decode_unit_io_macuio_0_bits_srcreq_5_idx),
    .io_macuio_0_bits_srcreq_5_busy(decode_unit_io_macuio_0_bits_srcreq_5_busy),
    .io_macuio_0_bits_srcreq_5_wkupidx_0(decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_0),
    .io_macuio_0_bits_srcreq_5_wkupidx_1(decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_1),
    .io_macuio_0_bits_srcreq_5_wkupidx_2(decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_2),
    .io_macuio_0_bits_srcreq_5_wkupidx_3(decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_3),
    .io_macuio_0_bits_srcreq_5_wkupidx_4(decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_4),
    .io_macuio_0_bits_srcreq_5_wkupidx_5(decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_5),
    .io_macuio_0_bits_wbvld(decode_unit_io_macuio_0_bits_wbvld),
    .io_macuio_0_bits_wbreq(decode_unit_io_macuio_0_bits_wbreq),
    .io_macuio_0_bits_waridx_0(decode_unit_io_macuio_0_bits_waridx_0),
    .io_macuio_0_bits_waridx_1(decode_unit_io_macuio_0_bits_waridx_1),
    .io_macuio_0_bits_waridx_2(decode_unit_io_macuio_0_bits_waridx_2),
    .io_macuio_0_bits_waridx_3(decode_unit_io_macuio_0_bits_waridx_3),
    .io_macuio_0_bits_waridx_4(decode_unit_io_macuio_0_bits_waridx_4),
    .io_macuio_0_bits_wawidx_0(decode_unit_io_macuio_0_bits_wawidx_0),
    .io_macuio_0_bits_wawidx_1(decode_unit_io_macuio_0_bits_wawidx_1),
    .io_macuio_0_bits_wawidx_2(decode_unit_io_macuio_0_bits_wawidx_2),
    .io_macuio_0_bits_wawidx_3(decode_unit_io_macuio_0_bits_wawidx_3),
    .io_macuio_0_bits_wawidx_4(decode_unit_io_macuio_0_bits_wawidx_4),
    .io_macuio_1_ready(decode_unit_io_macuio_1_ready),
    .io_macuio_1_valid(decode_unit_io_macuio_1_valid),
    .io_macuio_1_bits_vlen(decode_unit_io_macuio_1_bits_vlen),
    .io_macuio_1_bits_select(decode_unit_io_macuio_1_bits_select),
    .io_macuio_1_bits_drc(decode_unit_io_macuio_1_bits_drc),
    .io_macuio_1_bits_pow(decode_unit_io_macuio_1_bits_pow),
    .io_macuio_1_bits_loop(decode_unit_io_macuio_1_bits_loop),
    .io_macuio_1_bits_drcgain(decode_unit_io_macuio_1_bits_drcgain),
    .io_macuio_1_bits_drcnum(decode_unit_io_macuio_1_bits_drcnum),
    .io_macuio_1_bits_srcreq_0_valid(decode_unit_io_macuio_1_bits_srcreq_0_valid),
    .io_macuio_1_bits_srcreq_0_isgroup(decode_unit_io_macuio_1_bits_srcreq_0_isgroup),
    .io_macuio_1_bits_srcreq_0_iscoef(decode_unit_io_macuio_1_bits_srcreq_0_iscoef),
    .io_macuio_1_bits_srcreq_0_idx(decode_unit_io_macuio_1_bits_srcreq_0_idx),
    .io_macuio_1_bits_srcreq_0_busy(decode_unit_io_macuio_1_bits_srcreq_0_busy),
    .io_macuio_1_bits_srcreq_0_wkupidx_0(decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_0),
    .io_macuio_1_bits_srcreq_0_wkupidx_1(decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_1),
    .io_macuio_1_bits_srcreq_0_wkupidx_2(decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_2),
    .io_macuio_1_bits_srcreq_0_wkupidx_3(decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_3),
    .io_macuio_1_bits_srcreq_0_wkupidx_4(decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_4),
    .io_macuio_1_bits_srcreq_0_wkupidx_5(decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_5),
    .io_macuio_1_bits_srcreq_1_valid(decode_unit_io_macuio_1_bits_srcreq_1_valid),
    .io_macuio_1_bits_srcreq_1_isgroup(decode_unit_io_macuio_1_bits_srcreq_1_isgroup),
    .io_macuio_1_bits_srcreq_1_iscoef(decode_unit_io_macuio_1_bits_srcreq_1_iscoef),
    .io_macuio_1_bits_srcreq_1_idx(decode_unit_io_macuio_1_bits_srcreq_1_idx),
    .io_macuio_1_bits_srcreq_1_busy(decode_unit_io_macuio_1_bits_srcreq_1_busy),
    .io_macuio_1_bits_srcreq_1_wkupidx_0(decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_0),
    .io_macuio_1_bits_srcreq_1_wkupidx_1(decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_1),
    .io_macuio_1_bits_srcreq_1_wkupidx_2(decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_2),
    .io_macuio_1_bits_srcreq_1_wkupidx_3(decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_3),
    .io_macuio_1_bits_srcreq_1_wkupidx_4(decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_4),
    .io_macuio_1_bits_srcreq_1_wkupidx_5(decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_5),
    .io_macuio_1_bits_srcreq_2_valid(decode_unit_io_macuio_1_bits_srcreq_2_valid),
    .io_macuio_1_bits_srcreq_2_isgroup(decode_unit_io_macuio_1_bits_srcreq_2_isgroup),
    .io_macuio_1_bits_srcreq_2_iscoef(decode_unit_io_macuio_1_bits_srcreq_2_iscoef),
    .io_macuio_1_bits_srcreq_2_idx(decode_unit_io_macuio_1_bits_srcreq_2_idx),
    .io_macuio_1_bits_srcreq_2_busy(decode_unit_io_macuio_1_bits_srcreq_2_busy),
    .io_macuio_1_bits_srcreq_2_wkupidx_0(decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_0),
    .io_macuio_1_bits_srcreq_2_wkupidx_1(decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_1),
    .io_macuio_1_bits_srcreq_2_wkupidx_2(decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_2),
    .io_macuio_1_bits_srcreq_2_wkupidx_3(decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_3),
    .io_macuio_1_bits_srcreq_2_wkupidx_4(decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_4),
    .io_macuio_1_bits_srcreq_2_wkupidx_5(decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_5),
    .io_macuio_1_bits_srcreq_3_valid(decode_unit_io_macuio_1_bits_srcreq_3_valid),
    .io_macuio_1_bits_srcreq_3_isgroup(decode_unit_io_macuio_1_bits_srcreq_3_isgroup),
    .io_macuio_1_bits_srcreq_3_iscoef(decode_unit_io_macuio_1_bits_srcreq_3_iscoef),
    .io_macuio_1_bits_srcreq_3_idx(decode_unit_io_macuio_1_bits_srcreq_3_idx),
    .io_macuio_1_bits_srcreq_3_busy(decode_unit_io_macuio_1_bits_srcreq_3_busy),
    .io_macuio_1_bits_srcreq_3_wkupidx_0(decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_0),
    .io_macuio_1_bits_srcreq_3_wkupidx_1(decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_1),
    .io_macuio_1_bits_srcreq_3_wkupidx_2(decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_2),
    .io_macuio_1_bits_srcreq_3_wkupidx_3(decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_3),
    .io_macuio_1_bits_srcreq_3_wkupidx_4(decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_4),
    .io_macuio_1_bits_srcreq_3_wkupidx_5(decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_5),
    .io_macuio_1_bits_srcreq_4_valid(decode_unit_io_macuio_1_bits_srcreq_4_valid),
    .io_macuio_1_bits_srcreq_4_isgroup(decode_unit_io_macuio_1_bits_srcreq_4_isgroup),
    .io_macuio_1_bits_srcreq_4_iscoef(decode_unit_io_macuio_1_bits_srcreq_4_iscoef),
    .io_macuio_1_bits_srcreq_4_idx(decode_unit_io_macuio_1_bits_srcreq_4_idx),
    .io_macuio_1_bits_srcreq_4_busy(decode_unit_io_macuio_1_bits_srcreq_4_busy),
    .io_macuio_1_bits_srcreq_4_wkupidx_0(decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_0),
    .io_macuio_1_bits_srcreq_4_wkupidx_1(decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_1),
    .io_macuio_1_bits_srcreq_4_wkupidx_2(decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_2),
    .io_macuio_1_bits_srcreq_4_wkupidx_3(decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_3),
    .io_macuio_1_bits_srcreq_4_wkupidx_4(decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_4),
    .io_macuio_1_bits_srcreq_4_wkupidx_5(decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_5),
    .io_macuio_1_bits_srcreq_5_valid(decode_unit_io_macuio_1_bits_srcreq_5_valid),
    .io_macuio_1_bits_srcreq_5_isgroup(decode_unit_io_macuio_1_bits_srcreq_5_isgroup),
    .io_macuio_1_bits_srcreq_5_iscoef(decode_unit_io_macuio_1_bits_srcreq_5_iscoef),
    .io_macuio_1_bits_srcreq_5_idx(decode_unit_io_macuio_1_bits_srcreq_5_idx),
    .io_macuio_1_bits_srcreq_5_busy(decode_unit_io_macuio_1_bits_srcreq_5_busy),
    .io_macuio_1_bits_srcreq_5_wkupidx_0(decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_0),
    .io_macuio_1_bits_srcreq_5_wkupidx_1(decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_1),
    .io_macuio_1_bits_srcreq_5_wkupidx_2(decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_2),
    .io_macuio_1_bits_srcreq_5_wkupidx_3(decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_3),
    .io_macuio_1_bits_srcreq_5_wkupidx_4(decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_4),
    .io_macuio_1_bits_srcreq_5_wkupidx_5(decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_5),
    .io_macuio_1_bits_wbvld(decode_unit_io_macuio_1_bits_wbvld),
    .io_macuio_1_bits_wbreq(decode_unit_io_macuio_1_bits_wbreq),
    .io_macuio_1_bits_waridx_0(decode_unit_io_macuio_1_bits_waridx_0),
    .io_macuio_1_bits_waridx_1(decode_unit_io_macuio_1_bits_waridx_1),
    .io_macuio_1_bits_waridx_2(decode_unit_io_macuio_1_bits_waridx_2),
    .io_macuio_1_bits_waridx_3(decode_unit_io_macuio_1_bits_waridx_3),
    .io_macuio_1_bits_waridx_4(decode_unit_io_macuio_1_bits_waridx_4),
    .io_macuio_1_bits_wawidx_0(decode_unit_io_macuio_1_bits_wawidx_0),
    .io_macuio_1_bits_wawidx_1(decode_unit_io_macuio_1_bits_wawidx_1),
    .io_macuio_1_bits_wawidx_2(decode_unit_io_macuio_1_bits_wawidx_2),
    .io_macuio_1_bits_wawidx_3(decode_unit_io_macuio_1_bits_wawidx_3),
    .io_macuio_1_bits_wawidx_4(decode_unit_io_macuio_1_bits_wawidx_4),
    .io_macuio_2_ready(decode_unit_io_macuio_2_ready),
    .io_macuio_2_valid(decode_unit_io_macuio_2_valid),
    .io_macuio_2_bits_vlen(decode_unit_io_macuio_2_bits_vlen),
    .io_macuio_2_bits_select(decode_unit_io_macuio_2_bits_select),
    .io_macuio_2_bits_drc(decode_unit_io_macuio_2_bits_drc),
    .io_macuio_2_bits_pow(decode_unit_io_macuio_2_bits_pow),
    .io_macuio_2_bits_loop(decode_unit_io_macuio_2_bits_loop),
    .io_macuio_2_bits_drcgain(decode_unit_io_macuio_2_bits_drcgain),
    .io_macuio_2_bits_drcnum(decode_unit_io_macuio_2_bits_drcnum),
    .io_macuio_2_bits_srcreq_0_valid(decode_unit_io_macuio_2_bits_srcreq_0_valid),
    .io_macuio_2_bits_srcreq_0_isgroup(decode_unit_io_macuio_2_bits_srcreq_0_isgroup),
    .io_macuio_2_bits_srcreq_0_iscoef(decode_unit_io_macuio_2_bits_srcreq_0_iscoef),
    .io_macuio_2_bits_srcreq_0_idx(decode_unit_io_macuio_2_bits_srcreq_0_idx),
    .io_macuio_2_bits_srcreq_0_busy(decode_unit_io_macuio_2_bits_srcreq_0_busy),
    .io_macuio_2_bits_srcreq_0_wkupidx_0(decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_0),
    .io_macuio_2_bits_srcreq_0_wkupidx_1(decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_1),
    .io_macuio_2_bits_srcreq_0_wkupidx_2(decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_2),
    .io_macuio_2_bits_srcreq_0_wkupidx_3(decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_3),
    .io_macuio_2_bits_srcreq_0_wkupidx_4(decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_4),
    .io_macuio_2_bits_srcreq_0_wkupidx_5(decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_5),
    .io_macuio_2_bits_srcreq_1_valid(decode_unit_io_macuio_2_bits_srcreq_1_valid),
    .io_macuio_2_bits_srcreq_1_isgroup(decode_unit_io_macuio_2_bits_srcreq_1_isgroup),
    .io_macuio_2_bits_srcreq_1_iscoef(decode_unit_io_macuio_2_bits_srcreq_1_iscoef),
    .io_macuio_2_bits_srcreq_1_idx(decode_unit_io_macuio_2_bits_srcreq_1_idx),
    .io_macuio_2_bits_srcreq_1_busy(decode_unit_io_macuio_2_bits_srcreq_1_busy),
    .io_macuio_2_bits_srcreq_1_wkupidx_0(decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_0),
    .io_macuio_2_bits_srcreq_1_wkupidx_1(decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_1),
    .io_macuio_2_bits_srcreq_1_wkupidx_2(decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_2),
    .io_macuio_2_bits_srcreq_1_wkupidx_3(decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_3),
    .io_macuio_2_bits_srcreq_1_wkupidx_4(decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_4),
    .io_macuio_2_bits_srcreq_1_wkupidx_5(decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_5),
    .io_macuio_2_bits_srcreq_2_valid(decode_unit_io_macuio_2_bits_srcreq_2_valid),
    .io_macuio_2_bits_srcreq_2_isgroup(decode_unit_io_macuio_2_bits_srcreq_2_isgroup),
    .io_macuio_2_bits_srcreq_2_iscoef(decode_unit_io_macuio_2_bits_srcreq_2_iscoef),
    .io_macuio_2_bits_srcreq_2_idx(decode_unit_io_macuio_2_bits_srcreq_2_idx),
    .io_macuio_2_bits_srcreq_2_busy(decode_unit_io_macuio_2_bits_srcreq_2_busy),
    .io_macuio_2_bits_srcreq_2_wkupidx_0(decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_0),
    .io_macuio_2_bits_srcreq_2_wkupidx_1(decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_1),
    .io_macuio_2_bits_srcreq_2_wkupidx_2(decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_2),
    .io_macuio_2_bits_srcreq_2_wkupidx_3(decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_3),
    .io_macuio_2_bits_srcreq_2_wkupidx_4(decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_4),
    .io_macuio_2_bits_srcreq_2_wkupidx_5(decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_5),
    .io_macuio_2_bits_srcreq_3_valid(decode_unit_io_macuio_2_bits_srcreq_3_valid),
    .io_macuio_2_bits_srcreq_3_isgroup(decode_unit_io_macuio_2_bits_srcreq_3_isgroup),
    .io_macuio_2_bits_srcreq_3_iscoef(decode_unit_io_macuio_2_bits_srcreq_3_iscoef),
    .io_macuio_2_bits_srcreq_3_idx(decode_unit_io_macuio_2_bits_srcreq_3_idx),
    .io_macuio_2_bits_srcreq_3_busy(decode_unit_io_macuio_2_bits_srcreq_3_busy),
    .io_macuio_2_bits_srcreq_3_wkupidx_0(decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_0),
    .io_macuio_2_bits_srcreq_3_wkupidx_1(decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_1),
    .io_macuio_2_bits_srcreq_3_wkupidx_2(decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_2),
    .io_macuio_2_bits_srcreq_3_wkupidx_3(decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_3),
    .io_macuio_2_bits_srcreq_3_wkupidx_4(decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_4),
    .io_macuio_2_bits_srcreq_3_wkupidx_5(decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_5),
    .io_macuio_2_bits_srcreq_4_valid(decode_unit_io_macuio_2_bits_srcreq_4_valid),
    .io_macuio_2_bits_srcreq_4_isgroup(decode_unit_io_macuio_2_bits_srcreq_4_isgroup),
    .io_macuio_2_bits_srcreq_4_iscoef(decode_unit_io_macuio_2_bits_srcreq_4_iscoef),
    .io_macuio_2_bits_srcreq_4_idx(decode_unit_io_macuio_2_bits_srcreq_4_idx),
    .io_macuio_2_bits_srcreq_4_busy(decode_unit_io_macuio_2_bits_srcreq_4_busy),
    .io_macuio_2_bits_srcreq_4_wkupidx_0(decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_0),
    .io_macuio_2_bits_srcreq_4_wkupidx_1(decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_1),
    .io_macuio_2_bits_srcreq_4_wkupidx_2(decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_2),
    .io_macuio_2_bits_srcreq_4_wkupidx_3(decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_3),
    .io_macuio_2_bits_srcreq_4_wkupidx_4(decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_4),
    .io_macuio_2_bits_srcreq_4_wkupidx_5(decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_5),
    .io_macuio_2_bits_srcreq_5_valid(decode_unit_io_macuio_2_bits_srcreq_5_valid),
    .io_macuio_2_bits_srcreq_5_isgroup(decode_unit_io_macuio_2_bits_srcreq_5_isgroup),
    .io_macuio_2_bits_srcreq_5_iscoef(decode_unit_io_macuio_2_bits_srcreq_5_iscoef),
    .io_macuio_2_bits_srcreq_5_idx(decode_unit_io_macuio_2_bits_srcreq_5_idx),
    .io_macuio_2_bits_srcreq_5_busy(decode_unit_io_macuio_2_bits_srcreq_5_busy),
    .io_macuio_2_bits_srcreq_5_wkupidx_0(decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_0),
    .io_macuio_2_bits_srcreq_5_wkupidx_1(decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_1),
    .io_macuio_2_bits_srcreq_5_wkupidx_2(decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_2),
    .io_macuio_2_bits_srcreq_5_wkupidx_3(decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_3),
    .io_macuio_2_bits_srcreq_5_wkupidx_4(decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_4),
    .io_macuio_2_bits_srcreq_5_wkupidx_5(decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_5),
    .io_macuio_2_bits_wbvld(decode_unit_io_macuio_2_bits_wbvld),
    .io_macuio_2_bits_wbreq(decode_unit_io_macuio_2_bits_wbreq),
    .io_macuio_2_bits_waridx_0(decode_unit_io_macuio_2_bits_waridx_0),
    .io_macuio_2_bits_waridx_1(decode_unit_io_macuio_2_bits_waridx_1),
    .io_macuio_2_bits_waridx_2(decode_unit_io_macuio_2_bits_waridx_2),
    .io_macuio_2_bits_waridx_3(decode_unit_io_macuio_2_bits_waridx_3),
    .io_macuio_2_bits_waridx_4(decode_unit_io_macuio_2_bits_waridx_4),
    .io_macuio_2_bits_wawidx_0(decode_unit_io_macuio_2_bits_wawidx_0),
    .io_macuio_2_bits_wawidx_1(decode_unit_io_macuio_2_bits_wawidx_1),
    .io_macuio_2_bits_wawidx_2(decode_unit_io_macuio_2_bits_wawidx_2),
    .io_macuio_2_bits_wawidx_3(decode_unit_io_macuio_2_bits_wawidx_3),
    .io_macuio_2_bits_wawidx_4(decode_unit_io_macuio_2_bits_wawidx_4),
    .io_macuio_3_ready(decode_unit_io_macuio_3_ready),
    .io_macuio_3_valid(decode_unit_io_macuio_3_valid),
    .io_macuio_3_bits_vlen(decode_unit_io_macuio_3_bits_vlen),
    .io_macuio_3_bits_select(decode_unit_io_macuio_3_bits_select),
    .io_macuio_3_bits_drc(decode_unit_io_macuio_3_bits_drc),
    .io_macuio_3_bits_pow(decode_unit_io_macuio_3_bits_pow),
    .io_macuio_3_bits_loop(decode_unit_io_macuio_3_bits_loop),
    .io_macuio_3_bits_drcgain(decode_unit_io_macuio_3_bits_drcgain),
    .io_macuio_3_bits_drcnum(decode_unit_io_macuio_3_bits_drcnum),
    .io_macuio_3_bits_srcreq_0_valid(decode_unit_io_macuio_3_bits_srcreq_0_valid),
    .io_macuio_3_bits_srcreq_0_isgroup(decode_unit_io_macuio_3_bits_srcreq_0_isgroup),
    .io_macuio_3_bits_srcreq_0_iscoef(decode_unit_io_macuio_3_bits_srcreq_0_iscoef),
    .io_macuio_3_bits_srcreq_0_idx(decode_unit_io_macuio_3_bits_srcreq_0_idx),
    .io_macuio_3_bits_srcreq_0_busy(decode_unit_io_macuio_3_bits_srcreq_0_busy),
    .io_macuio_3_bits_srcreq_0_wkupidx_0(decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_0),
    .io_macuio_3_bits_srcreq_0_wkupidx_1(decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_1),
    .io_macuio_3_bits_srcreq_0_wkupidx_2(decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_2),
    .io_macuio_3_bits_srcreq_0_wkupidx_3(decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_3),
    .io_macuio_3_bits_srcreq_0_wkupidx_4(decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_4),
    .io_macuio_3_bits_srcreq_0_wkupidx_5(decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_5),
    .io_macuio_3_bits_srcreq_1_valid(decode_unit_io_macuio_3_bits_srcreq_1_valid),
    .io_macuio_3_bits_srcreq_1_isgroup(decode_unit_io_macuio_3_bits_srcreq_1_isgroup),
    .io_macuio_3_bits_srcreq_1_iscoef(decode_unit_io_macuio_3_bits_srcreq_1_iscoef),
    .io_macuio_3_bits_srcreq_1_idx(decode_unit_io_macuio_3_bits_srcreq_1_idx),
    .io_macuio_3_bits_srcreq_1_busy(decode_unit_io_macuio_3_bits_srcreq_1_busy),
    .io_macuio_3_bits_srcreq_1_wkupidx_0(decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_0),
    .io_macuio_3_bits_srcreq_1_wkupidx_1(decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_1),
    .io_macuio_3_bits_srcreq_1_wkupidx_2(decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_2),
    .io_macuio_3_bits_srcreq_1_wkupidx_3(decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_3),
    .io_macuio_3_bits_srcreq_1_wkupidx_4(decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_4),
    .io_macuio_3_bits_srcreq_1_wkupidx_5(decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_5),
    .io_macuio_3_bits_srcreq_2_valid(decode_unit_io_macuio_3_bits_srcreq_2_valid),
    .io_macuio_3_bits_srcreq_2_isgroup(decode_unit_io_macuio_3_bits_srcreq_2_isgroup),
    .io_macuio_3_bits_srcreq_2_iscoef(decode_unit_io_macuio_3_bits_srcreq_2_iscoef),
    .io_macuio_3_bits_srcreq_2_idx(decode_unit_io_macuio_3_bits_srcreq_2_idx),
    .io_macuio_3_bits_srcreq_2_busy(decode_unit_io_macuio_3_bits_srcreq_2_busy),
    .io_macuio_3_bits_srcreq_2_wkupidx_0(decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_0),
    .io_macuio_3_bits_srcreq_2_wkupidx_1(decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_1),
    .io_macuio_3_bits_srcreq_2_wkupidx_2(decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_2),
    .io_macuio_3_bits_srcreq_2_wkupidx_3(decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_3),
    .io_macuio_3_bits_srcreq_2_wkupidx_4(decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_4),
    .io_macuio_3_bits_srcreq_2_wkupidx_5(decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_5),
    .io_macuio_3_bits_srcreq_3_valid(decode_unit_io_macuio_3_bits_srcreq_3_valid),
    .io_macuio_3_bits_srcreq_3_isgroup(decode_unit_io_macuio_3_bits_srcreq_3_isgroup),
    .io_macuio_3_bits_srcreq_3_iscoef(decode_unit_io_macuio_3_bits_srcreq_3_iscoef),
    .io_macuio_3_bits_srcreq_3_idx(decode_unit_io_macuio_3_bits_srcreq_3_idx),
    .io_macuio_3_bits_srcreq_3_busy(decode_unit_io_macuio_3_bits_srcreq_3_busy),
    .io_macuio_3_bits_srcreq_3_wkupidx_0(decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_0),
    .io_macuio_3_bits_srcreq_3_wkupidx_1(decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_1),
    .io_macuio_3_bits_srcreq_3_wkupidx_2(decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_2),
    .io_macuio_3_bits_srcreq_3_wkupidx_3(decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_3),
    .io_macuio_3_bits_srcreq_3_wkupidx_4(decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_4),
    .io_macuio_3_bits_srcreq_3_wkupidx_5(decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_5),
    .io_macuio_3_bits_srcreq_4_valid(decode_unit_io_macuio_3_bits_srcreq_4_valid),
    .io_macuio_3_bits_srcreq_4_isgroup(decode_unit_io_macuio_3_bits_srcreq_4_isgroup),
    .io_macuio_3_bits_srcreq_4_iscoef(decode_unit_io_macuio_3_bits_srcreq_4_iscoef),
    .io_macuio_3_bits_srcreq_4_idx(decode_unit_io_macuio_3_bits_srcreq_4_idx),
    .io_macuio_3_bits_srcreq_4_busy(decode_unit_io_macuio_3_bits_srcreq_4_busy),
    .io_macuio_3_bits_srcreq_4_wkupidx_0(decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_0),
    .io_macuio_3_bits_srcreq_4_wkupidx_1(decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_1),
    .io_macuio_3_bits_srcreq_4_wkupidx_2(decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_2),
    .io_macuio_3_bits_srcreq_4_wkupidx_3(decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_3),
    .io_macuio_3_bits_srcreq_4_wkupidx_4(decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_4),
    .io_macuio_3_bits_srcreq_4_wkupidx_5(decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_5),
    .io_macuio_3_bits_srcreq_5_valid(decode_unit_io_macuio_3_bits_srcreq_5_valid),
    .io_macuio_3_bits_srcreq_5_isgroup(decode_unit_io_macuio_3_bits_srcreq_5_isgroup),
    .io_macuio_3_bits_srcreq_5_iscoef(decode_unit_io_macuio_3_bits_srcreq_5_iscoef),
    .io_macuio_3_bits_srcreq_5_idx(decode_unit_io_macuio_3_bits_srcreq_5_idx),
    .io_macuio_3_bits_srcreq_5_busy(decode_unit_io_macuio_3_bits_srcreq_5_busy),
    .io_macuio_3_bits_srcreq_5_wkupidx_0(decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_0),
    .io_macuio_3_bits_srcreq_5_wkupidx_1(decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_1),
    .io_macuio_3_bits_srcreq_5_wkupidx_2(decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_2),
    .io_macuio_3_bits_srcreq_5_wkupidx_3(decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_3),
    .io_macuio_3_bits_srcreq_5_wkupidx_4(decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_4),
    .io_macuio_3_bits_srcreq_5_wkupidx_5(decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_5),
    .io_macuio_3_bits_wbvld(decode_unit_io_macuio_3_bits_wbvld),
    .io_macuio_3_bits_wbreq(decode_unit_io_macuio_3_bits_wbreq),
    .io_macuio_3_bits_waridx_0(decode_unit_io_macuio_3_bits_waridx_0),
    .io_macuio_3_bits_waridx_1(decode_unit_io_macuio_3_bits_waridx_1),
    .io_macuio_3_bits_waridx_2(decode_unit_io_macuio_3_bits_waridx_2),
    .io_macuio_3_bits_waridx_3(decode_unit_io_macuio_3_bits_waridx_3),
    .io_macuio_3_bits_waridx_4(decode_unit_io_macuio_3_bits_waridx_4),
    .io_macuio_3_bits_wawidx_0(decode_unit_io_macuio_3_bits_wawidx_0),
    .io_macuio_3_bits_wawidx_1(decode_unit_io_macuio_3_bits_wawidx_1),
    .io_macuio_3_bits_wawidx_2(decode_unit_io_macuio_3_bits_wawidx_2),
    .io_macuio_3_bits_wawidx_3(decode_unit_io_macuio_3_bits_wawidx_3),
    .io_macuio_3_bits_wawidx_4(decode_unit_io_macuio_3_bits_wawidx_4),
    .io_macuio_4_ready(decode_unit_io_macuio_4_ready),
    .io_macuio_4_valid(decode_unit_io_macuio_4_valid),
    .io_macuio_4_bits_vlen(decode_unit_io_macuio_4_bits_vlen),
    .io_macuio_4_bits_select(decode_unit_io_macuio_4_bits_select),
    .io_macuio_4_bits_drc(decode_unit_io_macuio_4_bits_drc),
    .io_macuio_4_bits_pow(decode_unit_io_macuio_4_bits_pow),
    .io_macuio_4_bits_loop(decode_unit_io_macuio_4_bits_loop),
    .io_macuio_4_bits_drcgain(decode_unit_io_macuio_4_bits_drcgain),
    .io_macuio_4_bits_drcnum(decode_unit_io_macuio_4_bits_drcnum),
    .io_macuio_4_bits_srcreq_0_valid(decode_unit_io_macuio_4_bits_srcreq_0_valid),
    .io_macuio_4_bits_srcreq_0_isgroup(decode_unit_io_macuio_4_bits_srcreq_0_isgroup),
    .io_macuio_4_bits_srcreq_0_iscoef(decode_unit_io_macuio_4_bits_srcreq_0_iscoef),
    .io_macuio_4_bits_srcreq_0_idx(decode_unit_io_macuio_4_bits_srcreq_0_idx),
    .io_macuio_4_bits_srcreq_0_busy(decode_unit_io_macuio_4_bits_srcreq_0_busy),
    .io_macuio_4_bits_srcreq_0_wkupidx_0(decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_0),
    .io_macuio_4_bits_srcreq_0_wkupidx_1(decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_1),
    .io_macuio_4_bits_srcreq_0_wkupidx_2(decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_2),
    .io_macuio_4_bits_srcreq_0_wkupidx_3(decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_3),
    .io_macuio_4_bits_srcreq_0_wkupidx_4(decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_4),
    .io_macuio_4_bits_srcreq_0_wkupidx_5(decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_5),
    .io_macuio_4_bits_srcreq_1_valid(decode_unit_io_macuio_4_bits_srcreq_1_valid),
    .io_macuio_4_bits_srcreq_1_isgroup(decode_unit_io_macuio_4_bits_srcreq_1_isgroup),
    .io_macuio_4_bits_srcreq_1_iscoef(decode_unit_io_macuio_4_bits_srcreq_1_iscoef),
    .io_macuio_4_bits_srcreq_1_idx(decode_unit_io_macuio_4_bits_srcreq_1_idx),
    .io_macuio_4_bits_srcreq_1_busy(decode_unit_io_macuio_4_bits_srcreq_1_busy),
    .io_macuio_4_bits_srcreq_1_wkupidx_0(decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_0),
    .io_macuio_4_bits_srcreq_1_wkupidx_1(decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_1),
    .io_macuio_4_bits_srcreq_1_wkupidx_2(decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_2),
    .io_macuio_4_bits_srcreq_1_wkupidx_3(decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_3),
    .io_macuio_4_bits_srcreq_1_wkupidx_4(decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_4),
    .io_macuio_4_bits_srcreq_1_wkupidx_5(decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_5),
    .io_macuio_4_bits_srcreq_2_valid(decode_unit_io_macuio_4_bits_srcreq_2_valid),
    .io_macuio_4_bits_srcreq_2_isgroup(decode_unit_io_macuio_4_bits_srcreq_2_isgroup),
    .io_macuio_4_bits_srcreq_2_iscoef(decode_unit_io_macuio_4_bits_srcreq_2_iscoef),
    .io_macuio_4_bits_srcreq_2_idx(decode_unit_io_macuio_4_bits_srcreq_2_idx),
    .io_macuio_4_bits_srcreq_2_busy(decode_unit_io_macuio_4_bits_srcreq_2_busy),
    .io_macuio_4_bits_srcreq_2_wkupidx_0(decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_0),
    .io_macuio_4_bits_srcreq_2_wkupidx_1(decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_1),
    .io_macuio_4_bits_srcreq_2_wkupidx_2(decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_2),
    .io_macuio_4_bits_srcreq_2_wkupidx_3(decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_3),
    .io_macuio_4_bits_srcreq_2_wkupidx_4(decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_4),
    .io_macuio_4_bits_srcreq_2_wkupidx_5(decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_5),
    .io_macuio_4_bits_srcreq_3_valid(decode_unit_io_macuio_4_bits_srcreq_3_valid),
    .io_macuio_4_bits_srcreq_3_isgroup(decode_unit_io_macuio_4_bits_srcreq_3_isgroup),
    .io_macuio_4_bits_srcreq_3_iscoef(decode_unit_io_macuio_4_bits_srcreq_3_iscoef),
    .io_macuio_4_bits_srcreq_3_idx(decode_unit_io_macuio_4_bits_srcreq_3_idx),
    .io_macuio_4_bits_srcreq_3_busy(decode_unit_io_macuio_4_bits_srcreq_3_busy),
    .io_macuio_4_bits_srcreq_3_wkupidx_0(decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_0),
    .io_macuio_4_bits_srcreq_3_wkupidx_1(decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_1),
    .io_macuio_4_bits_srcreq_3_wkupidx_2(decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_2),
    .io_macuio_4_bits_srcreq_3_wkupidx_3(decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_3),
    .io_macuio_4_bits_srcreq_3_wkupidx_4(decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_4),
    .io_macuio_4_bits_srcreq_3_wkupidx_5(decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_5),
    .io_macuio_4_bits_srcreq_4_valid(decode_unit_io_macuio_4_bits_srcreq_4_valid),
    .io_macuio_4_bits_srcreq_4_isgroup(decode_unit_io_macuio_4_bits_srcreq_4_isgroup),
    .io_macuio_4_bits_srcreq_4_iscoef(decode_unit_io_macuio_4_bits_srcreq_4_iscoef),
    .io_macuio_4_bits_srcreq_4_idx(decode_unit_io_macuio_4_bits_srcreq_4_idx),
    .io_macuio_4_bits_srcreq_4_busy(decode_unit_io_macuio_4_bits_srcreq_4_busy),
    .io_macuio_4_bits_srcreq_4_wkupidx_0(decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_0),
    .io_macuio_4_bits_srcreq_4_wkupidx_1(decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_1),
    .io_macuio_4_bits_srcreq_4_wkupidx_2(decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_2),
    .io_macuio_4_bits_srcreq_4_wkupidx_3(decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_3),
    .io_macuio_4_bits_srcreq_4_wkupidx_4(decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_4),
    .io_macuio_4_bits_srcreq_4_wkupidx_5(decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_5),
    .io_macuio_4_bits_srcreq_5_valid(decode_unit_io_macuio_4_bits_srcreq_5_valid),
    .io_macuio_4_bits_srcreq_5_isgroup(decode_unit_io_macuio_4_bits_srcreq_5_isgroup),
    .io_macuio_4_bits_srcreq_5_iscoef(decode_unit_io_macuio_4_bits_srcreq_5_iscoef),
    .io_macuio_4_bits_srcreq_5_idx(decode_unit_io_macuio_4_bits_srcreq_5_idx),
    .io_macuio_4_bits_srcreq_5_busy(decode_unit_io_macuio_4_bits_srcreq_5_busy),
    .io_macuio_4_bits_srcreq_5_wkupidx_0(decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_0),
    .io_macuio_4_bits_srcreq_5_wkupidx_1(decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_1),
    .io_macuio_4_bits_srcreq_5_wkupidx_2(decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_2),
    .io_macuio_4_bits_srcreq_5_wkupidx_3(decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_3),
    .io_macuio_4_bits_srcreq_5_wkupidx_4(decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_4),
    .io_macuio_4_bits_srcreq_5_wkupidx_5(decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_5),
    .io_macuio_4_bits_wbvld(decode_unit_io_macuio_4_bits_wbvld),
    .io_macuio_4_bits_wbreq(decode_unit_io_macuio_4_bits_wbreq),
    .io_macuio_4_bits_waridx_0(decode_unit_io_macuio_4_bits_waridx_0),
    .io_macuio_4_bits_waridx_1(decode_unit_io_macuio_4_bits_waridx_1),
    .io_macuio_4_bits_waridx_2(decode_unit_io_macuio_4_bits_waridx_2),
    .io_macuio_4_bits_waridx_3(decode_unit_io_macuio_4_bits_waridx_3),
    .io_macuio_4_bits_waridx_4(decode_unit_io_macuio_4_bits_waridx_4),
    .io_macuio_4_bits_wawidx_0(decode_unit_io_macuio_4_bits_wawidx_0),
    .io_macuio_4_bits_wawidx_1(decode_unit_io_macuio_4_bits_wawidx_1),
    .io_macuio_4_bits_wawidx_2(decode_unit_io_macuio_4_bits_wawidx_2),
    .io_macuio_4_bits_wawidx_3(decode_unit_io_macuio_4_bits_wawidx_3),
    .io_macuio_4_bits_wawidx_4(decode_unit_io_macuio_4_bits_wawidx_4),
    .io_wd_check_0_valid(decode_unit_io_wd_check_0_valid),
    .io_wd_check_0_bits(decode_unit_io_wd_check_0_bits),
    .io_wd_check_1_valid(decode_unit_io_wd_check_1_valid),
    .io_wd_check_1_bits(decode_unit_io_wd_check_1_bits),
    .io_wd_check_2_valid(decode_unit_io_wd_check_2_valid),
    .io_wd_check_2_bits(decode_unit_io_wd_check_2_bits),
    .io_wd_check_3_valid(decode_unit_io_wd_check_3_valid),
    .io_wd_check_3_bits(decode_unit_io_wd_check_3_bits),
    .io_wd_check_4_valid(decode_unit_io_wd_check_4_valid),
    .io_wd_check_4_bits(decode_unit_io_wd_check_4_bits),
    .io_wd_check_5_valid(decode_unit_io_wd_check_5_valid),
    .io_wd_check_5_bits(decode_unit_io_wd_check_5_bits),
    .io_mac_r_check_0_0_valid(decode_unit_io_mac_r_check_0_0_valid),
    .io_mac_r_check_0_0_bits(decode_unit_io_mac_r_check_0_0_bits),
    .io_mac_r_check_0_1_valid(decode_unit_io_mac_r_check_0_1_valid),
    .io_mac_r_check_0_1_bits(decode_unit_io_mac_r_check_0_1_bits),
    .io_mac_r_check_0_2_valid(decode_unit_io_mac_r_check_0_2_valid),
    .io_mac_r_check_0_2_bits(decode_unit_io_mac_r_check_0_2_bits),
    .io_mac_r_check_0_3_valid(decode_unit_io_mac_r_check_0_3_valid),
    .io_mac_r_check_0_3_bits(decode_unit_io_mac_r_check_0_3_bits),
    .io_mac_r_check_0_4_valid(decode_unit_io_mac_r_check_0_4_valid),
    .io_mac_r_check_0_4_bits(decode_unit_io_mac_r_check_0_4_bits),
    .io_mac_r_check_0_5_valid(decode_unit_io_mac_r_check_0_5_valid),
    .io_mac_r_check_0_5_bits(decode_unit_io_mac_r_check_0_5_bits),
    .io_mac_r_check_1_0_valid(decode_unit_io_mac_r_check_1_0_valid),
    .io_mac_r_check_1_0_bits(decode_unit_io_mac_r_check_1_0_bits),
    .io_mac_r_check_1_1_valid(decode_unit_io_mac_r_check_1_1_valid),
    .io_mac_r_check_1_1_bits(decode_unit_io_mac_r_check_1_1_bits),
    .io_mac_r_check_1_2_valid(decode_unit_io_mac_r_check_1_2_valid),
    .io_mac_r_check_1_2_bits(decode_unit_io_mac_r_check_1_2_bits),
    .io_mac_r_check_1_3_valid(decode_unit_io_mac_r_check_1_3_valid),
    .io_mac_r_check_1_3_bits(decode_unit_io_mac_r_check_1_3_bits),
    .io_mac_r_check_1_4_valid(decode_unit_io_mac_r_check_1_4_valid),
    .io_mac_r_check_1_4_bits(decode_unit_io_mac_r_check_1_4_bits),
    .io_mac_r_check_1_5_valid(decode_unit_io_mac_r_check_1_5_valid),
    .io_mac_r_check_1_5_bits(decode_unit_io_mac_r_check_1_5_bits),
    .io_mac_r_check_2_0_valid(decode_unit_io_mac_r_check_2_0_valid),
    .io_mac_r_check_2_0_bits(decode_unit_io_mac_r_check_2_0_bits),
    .io_mac_r_check_2_1_valid(decode_unit_io_mac_r_check_2_1_valid),
    .io_mac_r_check_2_1_bits(decode_unit_io_mac_r_check_2_1_bits),
    .io_mac_r_check_2_2_valid(decode_unit_io_mac_r_check_2_2_valid),
    .io_mac_r_check_2_2_bits(decode_unit_io_mac_r_check_2_2_bits),
    .io_mac_r_check_2_3_valid(decode_unit_io_mac_r_check_2_3_valid),
    .io_mac_r_check_2_3_bits(decode_unit_io_mac_r_check_2_3_bits),
    .io_mac_r_check_2_4_valid(decode_unit_io_mac_r_check_2_4_valid),
    .io_mac_r_check_2_4_bits(decode_unit_io_mac_r_check_2_4_bits),
    .io_mac_r_check_2_5_valid(decode_unit_io_mac_r_check_2_5_valid),
    .io_mac_r_check_2_5_bits(decode_unit_io_mac_r_check_2_5_bits),
    .io_mac_r_check_3_0_valid(decode_unit_io_mac_r_check_3_0_valid),
    .io_mac_r_check_3_0_bits(decode_unit_io_mac_r_check_3_0_bits),
    .io_mac_r_check_3_1_valid(decode_unit_io_mac_r_check_3_1_valid),
    .io_mac_r_check_3_1_bits(decode_unit_io_mac_r_check_3_1_bits),
    .io_mac_r_check_3_2_valid(decode_unit_io_mac_r_check_3_2_valid),
    .io_mac_r_check_3_2_bits(decode_unit_io_mac_r_check_3_2_bits),
    .io_mac_r_check_3_3_valid(decode_unit_io_mac_r_check_3_3_valid),
    .io_mac_r_check_3_3_bits(decode_unit_io_mac_r_check_3_3_bits),
    .io_mac_r_check_3_4_valid(decode_unit_io_mac_r_check_3_4_valid),
    .io_mac_r_check_3_4_bits(decode_unit_io_mac_r_check_3_4_bits),
    .io_mac_r_check_3_5_valid(decode_unit_io_mac_r_check_3_5_valid),
    .io_mac_r_check_3_5_bits(decode_unit_io_mac_r_check_3_5_bits),
    .io_mac_r_check_4_0_valid(decode_unit_io_mac_r_check_4_0_valid),
    .io_mac_r_check_4_0_bits(decode_unit_io_mac_r_check_4_0_bits),
    .io_mac_r_check_4_1_valid(decode_unit_io_mac_r_check_4_1_valid),
    .io_mac_r_check_4_1_bits(decode_unit_io_mac_r_check_4_1_bits),
    .io_mac_r_check_4_2_valid(decode_unit_io_mac_r_check_4_2_valid),
    .io_mac_r_check_4_2_bits(decode_unit_io_mac_r_check_4_2_bits),
    .io_mac_r_check_4_3_valid(decode_unit_io_mac_r_check_4_3_valid),
    .io_mac_r_check_4_3_bits(decode_unit_io_mac_r_check_4_3_bits),
    .io_mac_r_check_4_4_valid(decode_unit_io_mac_r_check_4_4_valid),
    .io_mac_r_check_4_4_bits(decode_unit_io_mac_r_check_4_4_bits),
    .io_mac_r_check_4_5_valid(decode_unit_io_mac_r_check_4_5_valid),
    .io_mac_r_check_4_5_bits(decode_unit_io_mac_r_check_4_5_bits),
    .io_cor_r_check_0_valid(decode_unit_io_cor_r_check_0_valid),
    .io_cor_r_check_0_bits(decode_unit_io_cor_r_check_0_bits),
    .io_cor_r_check_1_valid(decode_unit_io_cor_r_check_1_valid),
    .io_cor_r_check_1_bits(decode_unit_io_cor_r_check_1_bits),
    .io_exuempty_0(decode_unit_io_exuempty_0),
    .io_exuempty_1(decode_unit_io_exuempty_1),
    .io_exuempty_2(decode_unit_io_exuempty_2),
    .io_exuempty_3(decode_unit_io_exuempty_3),
    .io_exuempty_4(decode_unit_io_exuempty_4),
    .io_exuempty_5(decode_unit_io_exuempty_5),
    .io_coruio_ready(decode_unit_io_coruio_ready),
    .io_coruio_valid(decode_unit_io_coruio_valid),
    .io_coruio_bits_cortype(decode_unit_io_coruio_bits_cortype),
    .io_coruio_bits_srcreq_0_valid(decode_unit_io_coruio_bits_srcreq_0_valid),
    .io_coruio_bits_srcreq_0_idx(decode_unit_io_coruio_bits_srcreq_0_idx),
    .io_coruio_bits_srcreq_0_busy(decode_unit_io_coruio_bits_srcreq_0_busy),
    .io_coruio_bits_srcreq_0_wkupidx_0(decode_unit_io_coruio_bits_srcreq_0_wkupidx_0),
    .io_coruio_bits_srcreq_0_wkupidx_1(decode_unit_io_coruio_bits_srcreq_0_wkupidx_1),
    .io_coruio_bits_srcreq_0_wkupidx_2(decode_unit_io_coruio_bits_srcreq_0_wkupidx_2),
    .io_coruio_bits_srcreq_0_wkupidx_3(decode_unit_io_coruio_bits_srcreq_0_wkupidx_3),
    .io_coruio_bits_srcreq_0_wkupidx_4(decode_unit_io_coruio_bits_srcreq_0_wkupidx_4),
    .io_coruio_bits_srcreq_0_wkupidx_5(decode_unit_io_coruio_bits_srcreq_0_wkupidx_5),
    .io_coruio_bits_srcreq_1_valid(decode_unit_io_coruio_bits_srcreq_1_valid),
    .io_coruio_bits_srcreq_1_idx(decode_unit_io_coruio_bits_srcreq_1_idx),
    .io_coruio_bits_srcreq_1_busy(decode_unit_io_coruio_bits_srcreq_1_busy),
    .io_coruio_bits_srcreq_1_wkupidx_0(decode_unit_io_coruio_bits_srcreq_1_wkupidx_0),
    .io_coruio_bits_srcreq_1_wkupidx_1(decode_unit_io_coruio_bits_srcreq_1_wkupidx_1),
    .io_coruio_bits_srcreq_1_wkupidx_2(decode_unit_io_coruio_bits_srcreq_1_wkupidx_2),
    .io_coruio_bits_srcreq_1_wkupidx_3(decode_unit_io_coruio_bits_srcreq_1_wkupidx_3),
    .io_coruio_bits_srcreq_1_wkupidx_4(decode_unit_io_coruio_bits_srcreq_1_wkupidx_4),
    .io_coruio_bits_srcreq_1_wkupidx_5(decode_unit_io_coruio_bits_srcreq_1_wkupidx_5),
    .io_coruio_bits_wbvld(decode_unit_io_coruio_bits_wbvld),
    .io_coruio_bits_wbreq(decode_unit_io_coruio_bits_wbreq),
    .io_coruio_bits_waridx_0(decode_unit_io_coruio_bits_waridx_0),
    .io_coruio_bits_waridx_1(decode_unit_io_coruio_bits_waridx_1),
    .io_coruio_bits_waridx_2(decode_unit_io_coruio_bits_waridx_2),
    .io_coruio_bits_waridx_3(decode_unit_io_coruio_bits_waridx_3),
    .io_coruio_bits_waridx_4(decode_unit_io_coruio_bits_waridx_4),
    .io_coruio_bits_wawidx_0(decode_unit_io_coruio_bits_wawidx_0),
    .io_coruio_bits_wawidx_1(decode_unit_io_coruio_bits_wawidx_1),
    .io_coruio_bits_wawidx_2(decode_unit_io_coruio_bits_wawidx_2),
    .io_coruio_bits_wawidx_3(decode_unit_io_coruio_bits_wawidx_3),
    .io_coruio_bits_wawidx_4(decode_unit_io_coruio_bits_wawidx_4),
    .io_writerf_valid(decode_unit_io_writerf_valid),
    .io_writerf_bits_0(decode_unit_io_writerf_bits_0),
    .io_writerf_bits_1(decode_unit_io_writerf_bits_1),
    .io_writerf_bits_2(decode_unit_io_writerf_bits_2),
    .io_writerf_bits_3(decode_unit_io_writerf_bits_3),
    .io_readrf_0(decode_unit_io_readrf_0),
    .io_readrf_1(decode_unit_io_readrf_1),
    .io_coef_in_mainch_ch0_inputsel(decode_unit_io_coef_in_mainch_ch0_inputsel),
    .io_coef_in_mainch_ch1_inputsel(decode_unit_io_coef_in_mainch_ch1_inputsel)
  );
  RegFile reg_file ( // @[dsptop.scala 87:27]
    .clock(reg_file_clock),
    .reset(reg_file_reset),
    .io_exe_rd_0_req_isgroup(reg_file_io_exe_rd_0_req_isgroup),
    .io_exe_rd_0_req_iscoef(reg_file_io_exe_rd_0_req_iscoef),
    .io_exe_rd_0_req_idx(reg_file_io_exe_rd_0_req_idx),
    .io_exe_rd_0_req_gidx(reg_file_io_exe_rd_0_req_gidx),
    .io_exe_rd_0_resp(reg_file_io_exe_rd_0_resp),
    .io_exe_rd_1_req_isgroup(reg_file_io_exe_rd_1_req_isgroup),
    .io_exe_rd_1_req_iscoef(reg_file_io_exe_rd_1_req_iscoef),
    .io_exe_rd_1_req_idx(reg_file_io_exe_rd_1_req_idx),
    .io_exe_rd_1_req_gidx(reg_file_io_exe_rd_1_req_gidx),
    .io_exe_rd_1_req_sel(reg_file_io_exe_rd_1_req_sel),
    .io_exe_rd_1_resp(reg_file_io_exe_rd_1_resp),
    .io_exe_rd_2_req_isgroup(reg_file_io_exe_rd_2_req_isgroup),
    .io_exe_rd_2_req_iscoef(reg_file_io_exe_rd_2_req_iscoef),
    .io_exe_rd_2_req_idx(reg_file_io_exe_rd_2_req_idx),
    .io_exe_rd_2_req_gidx(reg_file_io_exe_rd_2_req_gidx),
    .io_exe_rd_2_resp(reg_file_io_exe_rd_2_resp),
    .io_exe_rd_3_req_isgroup(reg_file_io_exe_rd_3_req_isgroup),
    .io_exe_rd_3_req_iscoef(reg_file_io_exe_rd_3_req_iscoef),
    .io_exe_rd_3_req_idx(reg_file_io_exe_rd_3_req_idx),
    .io_exe_rd_3_req_gidx(reg_file_io_exe_rd_3_req_gidx),
    .io_exe_rd_3_req_sel(reg_file_io_exe_rd_3_req_sel),
    .io_exe_rd_3_resp(reg_file_io_exe_rd_3_resp),
    .io_exe_rd_4_req_isgroup(reg_file_io_exe_rd_4_req_isgroup),
    .io_exe_rd_4_req_iscoef(reg_file_io_exe_rd_4_req_iscoef),
    .io_exe_rd_4_req_idx(reg_file_io_exe_rd_4_req_idx),
    .io_exe_rd_4_req_gidx(reg_file_io_exe_rd_4_req_gidx),
    .io_exe_rd_4_resp(reg_file_io_exe_rd_4_resp),
    .io_exe_rd_5_req_isgroup(reg_file_io_exe_rd_5_req_isgroup),
    .io_exe_rd_5_req_iscoef(reg_file_io_exe_rd_5_req_iscoef),
    .io_exe_rd_5_req_idx(reg_file_io_exe_rd_5_req_idx),
    .io_exe_rd_5_req_gidx(reg_file_io_exe_rd_5_req_gidx),
    .io_exe_rd_5_req_sel(reg_file_io_exe_rd_5_req_sel),
    .io_exe_rd_5_resp(reg_file_io_exe_rd_5_resp),
    .io_exe_rd_6_req_isgroup(reg_file_io_exe_rd_6_req_isgroup),
    .io_exe_rd_6_req_iscoef(reg_file_io_exe_rd_6_req_iscoef),
    .io_exe_rd_6_req_idx(reg_file_io_exe_rd_6_req_idx),
    .io_exe_rd_6_req_gidx(reg_file_io_exe_rd_6_req_gidx),
    .io_exe_rd_6_resp(reg_file_io_exe_rd_6_resp),
    .io_exe_rd_7_req_isgroup(reg_file_io_exe_rd_7_req_isgroup),
    .io_exe_rd_7_req_iscoef(reg_file_io_exe_rd_7_req_iscoef),
    .io_exe_rd_7_req_idx(reg_file_io_exe_rd_7_req_idx),
    .io_exe_rd_7_req_gidx(reg_file_io_exe_rd_7_req_gidx),
    .io_exe_rd_7_req_sel(reg_file_io_exe_rd_7_req_sel),
    .io_exe_rd_7_resp(reg_file_io_exe_rd_7_resp),
    .io_exe_rd_8_req_isgroup(reg_file_io_exe_rd_8_req_isgroup),
    .io_exe_rd_8_req_iscoef(reg_file_io_exe_rd_8_req_iscoef),
    .io_exe_rd_8_req_idx(reg_file_io_exe_rd_8_req_idx),
    .io_exe_rd_8_req_gidx(reg_file_io_exe_rd_8_req_gidx),
    .io_exe_rd_8_resp(reg_file_io_exe_rd_8_resp),
    .io_exe_rd_9_req_isgroup(reg_file_io_exe_rd_9_req_isgroup),
    .io_exe_rd_9_req_iscoef(reg_file_io_exe_rd_9_req_iscoef),
    .io_exe_rd_9_req_idx(reg_file_io_exe_rd_9_req_idx),
    .io_exe_rd_9_req_gidx(reg_file_io_exe_rd_9_req_gidx),
    .io_exe_rd_9_req_sel(reg_file_io_exe_rd_9_req_sel),
    .io_exe_rd_9_resp(reg_file_io_exe_rd_9_resp),
    .io_exe_rd_10_req_idx(reg_file_io_exe_rd_10_req_idx),
    .io_exe_rd_10_resp(reg_file_io_exe_rd_10_resp),
    .io_exe_rd_11_req_idx(reg_file_io_exe_rd_11_req_idx),
    .io_exe_rd_11_resp(reg_file_io_exe_rd_11_resp),
    .io_exe_wb_0_wdata1(reg_file_io_exe_wb_0_wdata1),
    .io_exe_wb_0_wdata2(reg_file_io_exe_wb_0_wdata2),
    .io_exe_wb_0_vld(reg_file_io_exe_wb_0_vld),
    .io_exe_wb_0_gregidx(reg_file_io_exe_wb_0_gregidx),
    .io_exe_wb_1_wdata1(reg_file_io_exe_wb_1_wdata1),
    .io_exe_wb_1_wdata2(reg_file_io_exe_wb_1_wdata2),
    .io_exe_wb_1_vld(reg_file_io_exe_wb_1_vld),
    .io_exe_wb_1_gregidx(reg_file_io_exe_wb_1_gregidx),
    .io_exe_wb_2_wdata1(reg_file_io_exe_wb_2_wdata1),
    .io_exe_wb_2_wdata2(reg_file_io_exe_wb_2_wdata2),
    .io_exe_wb_2_vld(reg_file_io_exe_wb_2_vld),
    .io_exe_wb_2_gregidx(reg_file_io_exe_wb_2_gregidx),
    .io_exe_wb_3_wdata1(reg_file_io_exe_wb_3_wdata1),
    .io_exe_wb_3_wdata2(reg_file_io_exe_wb_3_wdata2),
    .io_exe_wb_3_vld(reg_file_io_exe_wb_3_vld),
    .io_exe_wb_3_gregidx(reg_file_io_exe_wb_3_gregidx),
    .io_exe_wb_4_wdata1(reg_file_io_exe_wb_4_wdata1),
    .io_exe_wb_4_wdata2(reg_file_io_exe_wb_4_wdata2),
    .io_exe_wb_4_vld(reg_file_io_exe_wb_4_vld),
    .io_exe_wb_4_gregidx(reg_file_io_exe_wb_4_gregidx),
    .io_exe_wb_5_wdata2(reg_file_io_exe_wb_5_wdata2),
    .io_exe_wb_5_vld(reg_file_io_exe_wb_5_vld),
    .io_exe_wb_5_gregidx(reg_file_io_exe_wb_5_gregidx),
    .io_dec_wb_valid(reg_file_io_dec_wb_valid),
    .io_dec_wb_bits_0(reg_file_io_dec_wb_bits_0),
    .io_dec_wb_bits_1(reg_file_io_dec_wb_bits_1),
    .io_dec_wb_bits_2(reg_file_io_dec_wb_bits_2),
    .io_dec_wb_bits_3(reg_file_io_dec_wb_bits_3),
    .io_dec_rd_0(reg_file_io_dec_rd_0),
    .io_dec_rd_1(reg_file_io_dec_rd_1),
    .io_coef_in_subch_ch2mix_0(reg_file_io_coef_in_subch_ch2mix_0),
    .io_coef_in_subch_ch2mix_1(reg_file_io_coef_in_subch_ch2mix_1),
    .io_coef_in_subch_ch2mix_2(reg_file_io_coef_in_subch_ch2mix_2),
    .io_coef_in_subch_ch2bq_0_0(reg_file_io_coef_in_subch_ch2bq_0_0),
    .io_coef_in_subch_ch2bq_0_1(reg_file_io_coef_in_subch_ch2bq_0_1),
    .io_coef_in_subch_ch2bq_0_2(reg_file_io_coef_in_subch_ch2bq_0_2),
    .io_coef_in_subch_ch2bq_0_3(reg_file_io_coef_in_subch_ch2bq_0_3),
    .io_coef_in_subch_ch2bq_0_4(reg_file_io_coef_in_subch_ch2bq_0_4),
    .io_coef_in_subch_ch2vol(reg_file_io_coef_in_subch_ch2vol),
    .io_coef_in_subch_ch2volsel(reg_file_io_coef_in_subch_ch2volsel),
    .io_coef_in_subch_ch3sel(reg_file_io_coef_in_subch_ch3sel),
    .io_coef_in_subch_ch3mix_0(reg_file_io_coef_in_subch_ch3mix_0),
    .io_coef_in_subch_ch3mix_1(reg_file_io_coef_in_subch_ch3mix_1),
    .io_coef_in_subch_ch3bq_0_0(reg_file_io_coef_in_subch_ch3bq_0_0),
    .io_coef_in_subch_ch3bq_0_1(reg_file_io_coef_in_subch_ch3bq_0_1),
    .io_coef_in_subch_ch3bq_0_2(reg_file_io_coef_in_subch_ch3bq_0_2),
    .io_coef_in_subch_ch3bq_0_3(reg_file_io_coef_in_subch_ch3bq_0_3),
    .io_coef_in_subch_ch3bq_0_4(reg_file_io_coef_in_subch_ch3bq_0_4),
    .io_coef_in_subch_ch3bq_1_0(reg_file_io_coef_in_subch_ch3bq_1_0),
    .io_coef_in_subch_ch3bq_1_1(reg_file_io_coef_in_subch_ch3bq_1_1),
    .io_coef_in_subch_ch3bq_1_2(reg_file_io_coef_in_subch_ch3bq_1_2),
    .io_coef_in_subch_ch3bq_1_3(reg_file_io_coef_in_subch_ch3bq_1_3),
    .io_coef_in_subch_ch3bq_1_4(reg_file_io_coef_in_subch_ch3bq_1_4),
    .io_coef_in_subch_ch3vol(reg_file_io_coef_in_subch_ch3vol),
    .io_coef_in_subch_ch3volsel(reg_file_io_coef_in_subch_ch3volsel),
    .io_coef_in_subch_drc_pow_0(reg_file_io_coef_in_subch_drc_pow_0),
    .io_coef_in_subch_drc_pow_1(reg_file_io_coef_in_subch_drc_pow_1),
    .io_coef_in_subch_drc_smooth_0(reg_file_io_coef_in_subch_drc_smooth_0),
    .io_coef_in_subch_drc_smooth_1(reg_file_io_coef_in_subch_drc_smooth_1),
    .io_coef_in_subch_drc_smooth_2(reg_file_io_coef_in_subch_drc_smooth_2),
    .io_coef_in_subch_drc_smooth_3(reg_file_io_coef_in_subch_drc_smooth_3),
    .io_coef_in_subch_drc_ratio(reg_file_io_coef_in_subch_drc_ratio),
    .io_coef_in_mainch_ch0_bqcoef_0_0(reg_file_io_coef_in_mainch_ch0_bqcoef_0_0),
    .io_coef_in_mainch_ch0_bqcoef_0_1(reg_file_io_coef_in_mainch_ch0_bqcoef_0_1),
    .io_coef_in_mainch_ch0_bqcoef_0_2(reg_file_io_coef_in_mainch_ch0_bqcoef_0_2),
    .io_coef_in_mainch_ch0_bqcoef_0_3(reg_file_io_coef_in_mainch_ch0_bqcoef_0_3),
    .io_coef_in_mainch_ch0_bqcoef_0_4(reg_file_io_coef_in_mainch_ch0_bqcoef_0_4),
    .io_coef_in_mainch_ch0_bqcoef_1_0(reg_file_io_coef_in_mainch_ch0_bqcoef_1_0),
    .io_coef_in_mainch_ch0_bqcoef_1_1(reg_file_io_coef_in_mainch_ch0_bqcoef_1_1),
    .io_coef_in_mainch_ch0_bqcoef_1_2(reg_file_io_coef_in_mainch_ch0_bqcoef_1_2),
    .io_coef_in_mainch_ch0_bqcoef_1_3(reg_file_io_coef_in_mainch_ch0_bqcoef_1_3),
    .io_coef_in_mainch_ch0_bqcoef_1_4(reg_file_io_coef_in_mainch_ch0_bqcoef_1_4),
    .io_coef_in_mainch_ch0_bqcoef_2_0(reg_file_io_coef_in_mainch_ch0_bqcoef_2_0),
    .io_coef_in_mainch_ch0_bqcoef_2_1(reg_file_io_coef_in_mainch_ch0_bqcoef_2_1),
    .io_coef_in_mainch_ch0_bqcoef_2_2(reg_file_io_coef_in_mainch_ch0_bqcoef_2_2),
    .io_coef_in_mainch_ch0_bqcoef_2_3(reg_file_io_coef_in_mainch_ch0_bqcoef_2_3),
    .io_coef_in_mainch_ch0_bqcoef_2_4(reg_file_io_coef_in_mainch_ch0_bqcoef_2_4),
    .io_coef_in_mainch_ch0_bqcoef_3_0(reg_file_io_coef_in_mainch_ch0_bqcoef_3_0),
    .io_coef_in_mainch_ch0_bqcoef_3_1(reg_file_io_coef_in_mainch_ch0_bqcoef_3_1),
    .io_coef_in_mainch_ch0_bqcoef_3_2(reg_file_io_coef_in_mainch_ch0_bqcoef_3_2),
    .io_coef_in_mainch_ch0_bqcoef_3_3(reg_file_io_coef_in_mainch_ch0_bqcoef_3_3),
    .io_coef_in_mainch_ch0_bqcoef_3_4(reg_file_io_coef_in_mainch_ch0_bqcoef_3_4),
    .io_coef_in_mainch_ch0_bqcoef_4_0(reg_file_io_coef_in_mainch_ch0_bqcoef_4_0),
    .io_coef_in_mainch_ch0_bqcoef_4_1(reg_file_io_coef_in_mainch_ch0_bqcoef_4_1),
    .io_coef_in_mainch_ch0_bqcoef_4_2(reg_file_io_coef_in_mainch_ch0_bqcoef_4_2),
    .io_coef_in_mainch_ch0_bqcoef_4_3(reg_file_io_coef_in_mainch_ch0_bqcoef_4_3),
    .io_coef_in_mainch_ch0_bqcoef_4_4(reg_file_io_coef_in_mainch_ch0_bqcoef_4_4),
    .io_coef_in_mainch_ch0_bqcoef_5_0(reg_file_io_coef_in_mainch_ch0_bqcoef_5_0),
    .io_coef_in_mainch_ch0_bqcoef_5_1(reg_file_io_coef_in_mainch_ch0_bqcoef_5_1),
    .io_coef_in_mainch_ch0_bqcoef_5_2(reg_file_io_coef_in_mainch_ch0_bqcoef_5_2),
    .io_coef_in_mainch_ch0_bqcoef_5_3(reg_file_io_coef_in_mainch_ch0_bqcoef_5_3),
    .io_coef_in_mainch_ch0_bqcoef_5_4(reg_file_io_coef_in_mainch_ch0_bqcoef_5_4),
    .io_coef_in_mainch_ch0_bqcoef_6_0(reg_file_io_coef_in_mainch_ch0_bqcoef_6_0),
    .io_coef_in_mainch_ch0_bqcoef_6_1(reg_file_io_coef_in_mainch_ch0_bqcoef_6_1),
    .io_coef_in_mainch_ch0_bqcoef_6_2(reg_file_io_coef_in_mainch_ch0_bqcoef_6_2),
    .io_coef_in_mainch_ch0_bqcoef_6_3(reg_file_io_coef_in_mainch_ch0_bqcoef_6_3),
    .io_coef_in_mainch_ch0_bqcoef_6_4(reg_file_io_coef_in_mainch_ch0_bqcoef_6_4),
    .io_coef_in_mainch_ch0_bqcoef_7_0(reg_file_io_coef_in_mainch_ch0_bqcoef_7_0),
    .io_coef_in_mainch_ch0_bqcoef_7_1(reg_file_io_coef_in_mainch_ch0_bqcoef_7_1),
    .io_coef_in_mainch_ch0_bqcoef_7_2(reg_file_io_coef_in_mainch_ch0_bqcoef_7_2),
    .io_coef_in_mainch_ch0_bqcoef_7_3(reg_file_io_coef_in_mainch_ch0_bqcoef_7_3),
    .io_coef_in_mainch_ch0_bqcoef_7_4(reg_file_io_coef_in_mainch_ch0_bqcoef_7_4),
    .io_coef_in_mainch_ch0_bqcoef_8_0(reg_file_io_coef_in_mainch_ch0_bqcoef_8_0),
    .io_coef_in_mainch_ch0_bqcoef_8_1(reg_file_io_coef_in_mainch_ch0_bqcoef_8_1),
    .io_coef_in_mainch_ch0_bqcoef_8_2(reg_file_io_coef_in_mainch_ch0_bqcoef_8_2),
    .io_coef_in_mainch_ch0_bqcoef_8_3(reg_file_io_coef_in_mainch_ch0_bqcoef_8_3),
    .io_coef_in_mainch_ch0_bqcoef_8_4(reg_file_io_coef_in_mainch_ch0_bqcoef_8_4),
    .io_coef_in_mainch_ch0_inputmix_0_0(reg_file_io_coef_in_mainch_ch0_inputmix_0_0),
    .io_coef_in_mainch_ch0_inputmix_0_1(reg_file_io_coef_in_mainch_ch0_inputmix_0_1),
    .io_coef_in_mainch_ch0_inputmix_1_0(reg_file_io_coef_in_mainch_ch0_inputmix_1_0),
    .io_coef_in_mainch_ch0_inputmix_1_1(reg_file_io_coef_in_mainch_ch0_inputmix_1_1),
    .io_coef_in_mainch_ch0_vol(reg_file_io_coef_in_mainch_ch0_vol),
    .io_coef_in_mainch_ch0_outputmix_0(reg_file_io_coef_in_mainch_ch0_outputmix_0),
    .io_coef_in_mainch_ch0_outputmix_1(reg_file_io_coef_in_mainch_ch0_outputmix_1),
    .io_coef_in_mainch_ch0_outputmix_2(reg_file_io_coef_in_mainch_ch0_outputmix_2),
    .io_coef_in_mainch_ch0_prescale(reg_file_io_coef_in_mainch_ch0_prescale),
    .io_coef_in_mainch_ch0_postscale(reg_file_io_coef_in_mainch_ch0_postscale),
    .io_coef_in_mainch_ch1_bqcoef_0_0(reg_file_io_coef_in_mainch_ch1_bqcoef_0_0),
    .io_coef_in_mainch_ch1_bqcoef_0_1(reg_file_io_coef_in_mainch_ch1_bqcoef_0_1),
    .io_coef_in_mainch_ch1_bqcoef_0_2(reg_file_io_coef_in_mainch_ch1_bqcoef_0_2),
    .io_coef_in_mainch_ch1_bqcoef_0_3(reg_file_io_coef_in_mainch_ch1_bqcoef_0_3),
    .io_coef_in_mainch_ch1_bqcoef_0_4(reg_file_io_coef_in_mainch_ch1_bqcoef_0_4),
    .io_coef_in_mainch_ch1_bqcoef_1_0(reg_file_io_coef_in_mainch_ch1_bqcoef_1_0),
    .io_coef_in_mainch_ch1_bqcoef_1_1(reg_file_io_coef_in_mainch_ch1_bqcoef_1_1),
    .io_coef_in_mainch_ch1_bqcoef_1_2(reg_file_io_coef_in_mainch_ch1_bqcoef_1_2),
    .io_coef_in_mainch_ch1_bqcoef_1_3(reg_file_io_coef_in_mainch_ch1_bqcoef_1_3),
    .io_coef_in_mainch_ch1_bqcoef_1_4(reg_file_io_coef_in_mainch_ch1_bqcoef_1_4),
    .io_coef_in_mainch_ch1_bqcoef_2_0(reg_file_io_coef_in_mainch_ch1_bqcoef_2_0),
    .io_coef_in_mainch_ch1_bqcoef_2_1(reg_file_io_coef_in_mainch_ch1_bqcoef_2_1),
    .io_coef_in_mainch_ch1_bqcoef_2_2(reg_file_io_coef_in_mainch_ch1_bqcoef_2_2),
    .io_coef_in_mainch_ch1_bqcoef_2_3(reg_file_io_coef_in_mainch_ch1_bqcoef_2_3),
    .io_coef_in_mainch_ch1_bqcoef_2_4(reg_file_io_coef_in_mainch_ch1_bqcoef_2_4),
    .io_coef_in_mainch_ch1_bqcoef_3_0(reg_file_io_coef_in_mainch_ch1_bqcoef_3_0),
    .io_coef_in_mainch_ch1_bqcoef_3_1(reg_file_io_coef_in_mainch_ch1_bqcoef_3_1),
    .io_coef_in_mainch_ch1_bqcoef_3_2(reg_file_io_coef_in_mainch_ch1_bqcoef_3_2),
    .io_coef_in_mainch_ch1_bqcoef_3_3(reg_file_io_coef_in_mainch_ch1_bqcoef_3_3),
    .io_coef_in_mainch_ch1_bqcoef_3_4(reg_file_io_coef_in_mainch_ch1_bqcoef_3_4),
    .io_coef_in_mainch_ch1_bqcoef_4_0(reg_file_io_coef_in_mainch_ch1_bqcoef_4_0),
    .io_coef_in_mainch_ch1_bqcoef_4_1(reg_file_io_coef_in_mainch_ch1_bqcoef_4_1),
    .io_coef_in_mainch_ch1_bqcoef_4_2(reg_file_io_coef_in_mainch_ch1_bqcoef_4_2),
    .io_coef_in_mainch_ch1_bqcoef_4_3(reg_file_io_coef_in_mainch_ch1_bqcoef_4_3),
    .io_coef_in_mainch_ch1_bqcoef_4_4(reg_file_io_coef_in_mainch_ch1_bqcoef_4_4),
    .io_coef_in_mainch_ch1_bqcoef_5_0(reg_file_io_coef_in_mainch_ch1_bqcoef_5_0),
    .io_coef_in_mainch_ch1_bqcoef_5_1(reg_file_io_coef_in_mainch_ch1_bqcoef_5_1),
    .io_coef_in_mainch_ch1_bqcoef_5_2(reg_file_io_coef_in_mainch_ch1_bqcoef_5_2),
    .io_coef_in_mainch_ch1_bqcoef_5_3(reg_file_io_coef_in_mainch_ch1_bqcoef_5_3),
    .io_coef_in_mainch_ch1_bqcoef_5_4(reg_file_io_coef_in_mainch_ch1_bqcoef_5_4),
    .io_coef_in_mainch_ch1_bqcoef_6_0(reg_file_io_coef_in_mainch_ch1_bqcoef_6_0),
    .io_coef_in_mainch_ch1_bqcoef_6_1(reg_file_io_coef_in_mainch_ch1_bqcoef_6_1),
    .io_coef_in_mainch_ch1_bqcoef_6_2(reg_file_io_coef_in_mainch_ch1_bqcoef_6_2),
    .io_coef_in_mainch_ch1_bqcoef_6_3(reg_file_io_coef_in_mainch_ch1_bqcoef_6_3),
    .io_coef_in_mainch_ch1_bqcoef_6_4(reg_file_io_coef_in_mainch_ch1_bqcoef_6_4),
    .io_coef_in_mainch_ch1_bqcoef_7_0(reg_file_io_coef_in_mainch_ch1_bqcoef_7_0),
    .io_coef_in_mainch_ch1_bqcoef_7_1(reg_file_io_coef_in_mainch_ch1_bqcoef_7_1),
    .io_coef_in_mainch_ch1_bqcoef_7_2(reg_file_io_coef_in_mainch_ch1_bqcoef_7_2),
    .io_coef_in_mainch_ch1_bqcoef_7_3(reg_file_io_coef_in_mainch_ch1_bqcoef_7_3),
    .io_coef_in_mainch_ch1_bqcoef_7_4(reg_file_io_coef_in_mainch_ch1_bqcoef_7_4),
    .io_coef_in_mainch_ch1_bqcoef_8_0(reg_file_io_coef_in_mainch_ch1_bqcoef_8_0),
    .io_coef_in_mainch_ch1_bqcoef_8_1(reg_file_io_coef_in_mainch_ch1_bqcoef_8_1),
    .io_coef_in_mainch_ch1_bqcoef_8_2(reg_file_io_coef_in_mainch_ch1_bqcoef_8_2),
    .io_coef_in_mainch_ch1_bqcoef_8_3(reg_file_io_coef_in_mainch_ch1_bqcoef_8_3),
    .io_coef_in_mainch_ch1_bqcoef_8_4(reg_file_io_coef_in_mainch_ch1_bqcoef_8_4),
    .io_coef_in_mainch_ch1_inputmix_0_0(reg_file_io_coef_in_mainch_ch1_inputmix_0_0),
    .io_coef_in_mainch_ch1_inputmix_0_1(reg_file_io_coef_in_mainch_ch1_inputmix_0_1),
    .io_coef_in_mainch_ch1_inputmix_1_0(reg_file_io_coef_in_mainch_ch1_inputmix_1_0),
    .io_coef_in_mainch_ch1_inputmix_1_1(reg_file_io_coef_in_mainch_ch1_inputmix_1_1),
    .io_coef_in_mainch_ch1_vol(reg_file_io_coef_in_mainch_ch1_vol),
    .io_coef_in_mainch_ch1_outputmix_0(reg_file_io_coef_in_mainch_ch1_outputmix_0),
    .io_coef_in_mainch_ch1_outputmix_1(reg_file_io_coef_in_mainch_ch1_outputmix_1),
    .io_coef_in_mainch_ch1_outputmix_2(reg_file_io_coef_in_mainch_ch1_outputmix_2),
    .io_coef_in_mainch_drc_pow_0(reg_file_io_coef_in_mainch_drc_pow_0),
    .io_coef_in_mainch_drc_pow_1(reg_file_io_coef_in_mainch_drc_pow_1),
    .io_coef_in_mainch_drc_smooth_0(reg_file_io_coef_in_mainch_drc_smooth_0),
    .io_coef_in_mainch_drc_smooth_1(reg_file_io_coef_in_mainch_drc_smooth_1),
    .io_coef_in_mainch_drc_smooth_2(reg_file_io_coef_in_mainch_drc_smooth_2),
    .io_coef_in_mainch_drc_smooth_3(reg_file_io_coef_in_mainch_drc_smooth_3),
    .io_coef_in_mainch_drc_ratio(reg_file_io_coef_in_mainch_drc_ratio)
  );
  MacUnit mac_units_0 ( // @[dsptop.scala 88:70]
    .clock(mac_units_0_clock),
    .reset(mac_units_0_reset),
    .io_uopin_ready(mac_units_0_io_uopin_ready),
    .io_uopin_valid(mac_units_0_io_uopin_valid),
    .io_uopin_bits_vlen(mac_units_0_io_uopin_bits_vlen),
    .io_uopin_bits_select(mac_units_0_io_uopin_bits_select),
    .io_uopin_bits_drc(mac_units_0_io_uopin_bits_drc),
    .io_uopin_bits_pow(mac_units_0_io_uopin_bits_pow),
    .io_uopin_bits_loop(mac_units_0_io_uopin_bits_loop),
    .io_uopin_bits_drcgain(mac_units_0_io_uopin_bits_drcgain),
    .io_uopin_bits_drcnum(mac_units_0_io_uopin_bits_drcnum),
    .io_uopin_bits_srcreq_0_valid(mac_units_0_io_uopin_bits_srcreq_0_valid),
    .io_uopin_bits_srcreq_0_isgroup(mac_units_0_io_uopin_bits_srcreq_0_isgroup),
    .io_uopin_bits_srcreq_0_iscoef(mac_units_0_io_uopin_bits_srcreq_0_iscoef),
    .io_uopin_bits_srcreq_0_idx(mac_units_0_io_uopin_bits_srcreq_0_idx),
    .io_uopin_bits_srcreq_0_busy(mac_units_0_io_uopin_bits_srcreq_0_busy),
    .io_uopin_bits_srcreq_0_wkupidx_0(mac_units_0_io_uopin_bits_srcreq_0_wkupidx_0),
    .io_uopin_bits_srcreq_0_wkupidx_1(mac_units_0_io_uopin_bits_srcreq_0_wkupidx_1),
    .io_uopin_bits_srcreq_0_wkupidx_2(mac_units_0_io_uopin_bits_srcreq_0_wkupidx_2),
    .io_uopin_bits_srcreq_0_wkupidx_3(mac_units_0_io_uopin_bits_srcreq_0_wkupidx_3),
    .io_uopin_bits_srcreq_0_wkupidx_4(mac_units_0_io_uopin_bits_srcreq_0_wkupidx_4),
    .io_uopin_bits_srcreq_0_wkupidx_5(mac_units_0_io_uopin_bits_srcreq_0_wkupidx_5),
    .io_uopin_bits_srcreq_1_valid(mac_units_0_io_uopin_bits_srcreq_1_valid),
    .io_uopin_bits_srcreq_1_isgroup(mac_units_0_io_uopin_bits_srcreq_1_isgroup),
    .io_uopin_bits_srcreq_1_iscoef(mac_units_0_io_uopin_bits_srcreq_1_iscoef),
    .io_uopin_bits_srcreq_1_idx(mac_units_0_io_uopin_bits_srcreq_1_idx),
    .io_uopin_bits_srcreq_1_busy(mac_units_0_io_uopin_bits_srcreq_1_busy),
    .io_uopin_bits_srcreq_1_wkupidx_0(mac_units_0_io_uopin_bits_srcreq_1_wkupidx_0),
    .io_uopin_bits_srcreq_1_wkupidx_1(mac_units_0_io_uopin_bits_srcreq_1_wkupidx_1),
    .io_uopin_bits_srcreq_1_wkupidx_2(mac_units_0_io_uopin_bits_srcreq_1_wkupidx_2),
    .io_uopin_bits_srcreq_1_wkupidx_3(mac_units_0_io_uopin_bits_srcreq_1_wkupidx_3),
    .io_uopin_bits_srcreq_1_wkupidx_4(mac_units_0_io_uopin_bits_srcreq_1_wkupidx_4),
    .io_uopin_bits_srcreq_1_wkupidx_5(mac_units_0_io_uopin_bits_srcreq_1_wkupidx_5),
    .io_uopin_bits_srcreq_2_valid(mac_units_0_io_uopin_bits_srcreq_2_valid),
    .io_uopin_bits_srcreq_2_isgroup(mac_units_0_io_uopin_bits_srcreq_2_isgroup),
    .io_uopin_bits_srcreq_2_iscoef(mac_units_0_io_uopin_bits_srcreq_2_iscoef),
    .io_uopin_bits_srcreq_2_idx(mac_units_0_io_uopin_bits_srcreq_2_idx),
    .io_uopin_bits_srcreq_2_busy(mac_units_0_io_uopin_bits_srcreq_2_busy),
    .io_uopin_bits_srcreq_2_wkupidx_0(mac_units_0_io_uopin_bits_srcreq_2_wkupidx_0),
    .io_uopin_bits_srcreq_2_wkupidx_1(mac_units_0_io_uopin_bits_srcreq_2_wkupidx_1),
    .io_uopin_bits_srcreq_2_wkupidx_2(mac_units_0_io_uopin_bits_srcreq_2_wkupidx_2),
    .io_uopin_bits_srcreq_2_wkupidx_3(mac_units_0_io_uopin_bits_srcreq_2_wkupidx_3),
    .io_uopin_bits_srcreq_2_wkupidx_4(mac_units_0_io_uopin_bits_srcreq_2_wkupidx_4),
    .io_uopin_bits_srcreq_2_wkupidx_5(mac_units_0_io_uopin_bits_srcreq_2_wkupidx_5),
    .io_uopin_bits_srcreq_3_valid(mac_units_0_io_uopin_bits_srcreq_3_valid),
    .io_uopin_bits_srcreq_3_isgroup(mac_units_0_io_uopin_bits_srcreq_3_isgroup),
    .io_uopin_bits_srcreq_3_iscoef(mac_units_0_io_uopin_bits_srcreq_3_iscoef),
    .io_uopin_bits_srcreq_3_idx(mac_units_0_io_uopin_bits_srcreq_3_idx),
    .io_uopin_bits_srcreq_3_busy(mac_units_0_io_uopin_bits_srcreq_3_busy),
    .io_uopin_bits_srcreq_3_wkupidx_0(mac_units_0_io_uopin_bits_srcreq_3_wkupidx_0),
    .io_uopin_bits_srcreq_3_wkupidx_1(mac_units_0_io_uopin_bits_srcreq_3_wkupidx_1),
    .io_uopin_bits_srcreq_3_wkupidx_2(mac_units_0_io_uopin_bits_srcreq_3_wkupidx_2),
    .io_uopin_bits_srcreq_3_wkupidx_3(mac_units_0_io_uopin_bits_srcreq_3_wkupidx_3),
    .io_uopin_bits_srcreq_3_wkupidx_4(mac_units_0_io_uopin_bits_srcreq_3_wkupidx_4),
    .io_uopin_bits_srcreq_3_wkupidx_5(mac_units_0_io_uopin_bits_srcreq_3_wkupidx_5),
    .io_uopin_bits_srcreq_4_valid(mac_units_0_io_uopin_bits_srcreq_4_valid),
    .io_uopin_bits_srcreq_4_isgroup(mac_units_0_io_uopin_bits_srcreq_4_isgroup),
    .io_uopin_bits_srcreq_4_iscoef(mac_units_0_io_uopin_bits_srcreq_4_iscoef),
    .io_uopin_bits_srcreq_4_idx(mac_units_0_io_uopin_bits_srcreq_4_idx),
    .io_uopin_bits_srcreq_4_busy(mac_units_0_io_uopin_bits_srcreq_4_busy),
    .io_uopin_bits_srcreq_4_wkupidx_0(mac_units_0_io_uopin_bits_srcreq_4_wkupidx_0),
    .io_uopin_bits_srcreq_4_wkupidx_1(mac_units_0_io_uopin_bits_srcreq_4_wkupidx_1),
    .io_uopin_bits_srcreq_4_wkupidx_2(mac_units_0_io_uopin_bits_srcreq_4_wkupidx_2),
    .io_uopin_bits_srcreq_4_wkupidx_3(mac_units_0_io_uopin_bits_srcreq_4_wkupidx_3),
    .io_uopin_bits_srcreq_4_wkupidx_4(mac_units_0_io_uopin_bits_srcreq_4_wkupidx_4),
    .io_uopin_bits_srcreq_4_wkupidx_5(mac_units_0_io_uopin_bits_srcreq_4_wkupidx_5),
    .io_uopin_bits_srcreq_5_valid(mac_units_0_io_uopin_bits_srcreq_5_valid),
    .io_uopin_bits_srcreq_5_isgroup(mac_units_0_io_uopin_bits_srcreq_5_isgroup),
    .io_uopin_bits_srcreq_5_iscoef(mac_units_0_io_uopin_bits_srcreq_5_iscoef),
    .io_uopin_bits_srcreq_5_idx(mac_units_0_io_uopin_bits_srcreq_5_idx),
    .io_uopin_bits_srcreq_5_busy(mac_units_0_io_uopin_bits_srcreq_5_busy),
    .io_uopin_bits_srcreq_5_wkupidx_0(mac_units_0_io_uopin_bits_srcreq_5_wkupidx_0),
    .io_uopin_bits_srcreq_5_wkupidx_1(mac_units_0_io_uopin_bits_srcreq_5_wkupidx_1),
    .io_uopin_bits_srcreq_5_wkupidx_2(mac_units_0_io_uopin_bits_srcreq_5_wkupidx_2),
    .io_uopin_bits_srcreq_5_wkupidx_3(mac_units_0_io_uopin_bits_srcreq_5_wkupidx_3),
    .io_uopin_bits_srcreq_5_wkupidx_4(mac_units_0_io_uopin_bits_srcreq_5_wkupidx_4),
    .io_uopin_bits_srcreq_5_wkupidx_5(mac_units_0_io_uopin_bits_srcreq_5_wkupidx_5),
    .io_uopin_bits_wbvld(mac_units_0_io_uopin_bits_wbvld),
    .io_uopin_bits_wbreq(mac_units_0_io_uopin_bits_wbreq),
    .io_uopin_bits_waridx_0(mac_units_0_io_uopin_bits_waridx_0),
    .io_uopin_bits_waridx_1(mac_units_0_io_uopin_bits_waridx_1),
    .io_uopin_bits_waridx_2(mac_units_0_io_uopin_bits_waridx_2),
    .io_uopin_bits_waridx_3(mac_units_0_io_uopin_bits_waridx_3),
    .io_uopin_bits_waridx_4(mac_units_0_io_uopin_bits_waridx_4),
    .io_uopin_bits_wawidx_0(mac_units_0_io_uopin_bits_wawidx_0),
    .io_uopin_bits_wawidx_1(mac_units_0_io_uopin_bits_wawidx_1),
    .io_uopin_bits_wawidx_2(mac_units_0_io_uopin_bits_wawidx_2),
    .io_uopin_bits_wawidx_3(mac_units_0_io_uopin_bits_wawidx_3),
    .io_uopin_bits_wawidx_4(mac_units_0_io_uopin_bits_wawidx_4),
    .io_rfreq_0_req_isgroup(mac_units_0_io_rfreq_0_req_isgroup),
    .io_rfreq_0_req_iscoef(mac_units_0_io_rfreq_0_req_iscoef),
    .io_rfreq_0_req_idx(mac_units_0_io_rfreq_0_req_idx),
    .io_rfreq_0_req_gidx(mac_units_0_io_rfreq_0_req_gidx),
    .io_rfreq_0_resp(mac_units_0_io_rfreq_0_resp),
    .io_rfreq_1_req_isgroup(mac_units_0_io_rfreq_1_req_isgroup),
    .io_rfreq_1_req_iscoef(mac_units_0_io_rfreq_1_req_iscoef),
    .io_rfreq_1_req_idx(mac_units_0_io_rfreq_1_req_idx),
    .io_rfreq_1_req_gidx(mac_units_0_io_rfreq_1_req_gidx),
    .io_rfreq_1_req_sel(mac_units_0_io_rfreq_1_req_sel),
    .io_rfreq_1_resp(mac_units_0_io_rfreq_1_resp),
    .io_wbreq_wdata1(mac_units_0_io_wbreq_wdata1),
    .io_wbreq_wdata2(mac_units_0_io_wbreq_wdata2),
    .io_wbreq_vld(mac_units_0_io_wbreq_vld),
    .io_wbreq_gregidx(mac_units_0_io_wbreq_gregidx),
    .io_fwd_wkup_valid(mac_units_0_io_fwd_wkup_valid),
    .io_fwd_wkup_bits(mac_units_0_io_fwd_wkup_bits),
    .io_empty(mac_units_0_io_empty),
    .io_raw_wkup_0_valid(mac_units_0_io_raw_wkup_0_valid),
    .io_raw_wkup_0_bits(mac_units_0_io_raw_wkup_0_bits),
    .io_raw_wkup_1_valid(mac_units_0_io_raw_wkup_1_valid),
    .io_raw_wkup_1_bits(mac_units_0_io_raw_wkup_1_bits),
    .io_raw_wkup_2_valid(mac_units_0_io_raw_wkup_2_valid),
    .io_raw_wkup_2_bits(mac_units_0_io_raw_wkup_2_bits),
    .io_raw_wkup_3_valid(mac_units_0_io_raw_wkup_3_valid),
    .io_raw_wkup_3_bits(mac_units_0_io_raw_wkup_3_bits),
    .io_raw_wkup_4_valid(mac_units_0_io_raw_wkup_4_valid),
    .io_raw_wkup_4_bits(mac_units_0_io_raw_wkup_4_bits),
    .io_raw_wkup_5_valid(mac_units_0_io_raw_wkup_5_valid),
    .io_raw_wkup_5_bits(mac_units_0_io_raw_wkup_5_bits),
    .io_wbcheck_valid(mac_units_0_io_wbcheck_valid),
    .io_wbcheck_bits(mac_units_0_io_wbcheck_bits),
    .io_r_check_0_valid(mac_units_0_io_r_check_0_valid),
    .io_r_check_0_bits(mac_units_0_io_r_check_0_bits),
    .io_r_check_1_valid(mac_units_0_io_r_check_1_valid),
    .io_r_check_1_bits(mac_units_0_io_r_check_1_bits),
    .io_r_check_2_valid(mac_units_0_io_r_check_2_valid),
    .io_r_check_2_bits(mac_units_0_io_r_check_2_bits),
    .io_r_check_3_valid(mac_units_0_io_r_check_3_valid),
    .io_r_check_3_bits(mac_units_0_io_r_check_3_bits),
    .io_r_check_4_valid(mac_units_0_io_r_check_4_valid),
    .io_r_check_4_bits(mac_units_0_io_r_check_4_bits),
    .io_r_check_5_valid(mac_units_0_io_r_check_5_valid),
    .io_r_check_5_bits(mac_units_0_io_r_check_5_bits),
    .io_other_flop_0(mac_units_0_io_other_flop_0),
    .io_other_flop_1(mac_units_0_io_other_flop_1),
    .io_other_flop_2(mac_units_0_io_other_flop_2),
    .io_other_flop_3(mac_units_0_io_other_flop_3),
    .io_other_flop_4(mac_units_0_io_other_flop_4),
    .io_flop(mac_units_0_io_flop),
    .io_coef_subch_drc_th(mac_units_0_io_coef_subch_drc_th),
    .io_coef_subch_drc_offset(mac_units_0_io_coef_subch_drc_offset),
    .io_coef_subch_drc_drcen(mac_units_0_io_coef_subch_drc_drcen),
    .io_coef_mainch_ch0_autoloop(mac_units_0_io_coef_mainch_ch0_autoloop),
    .io_coef_mainch_drc_th(mac_units_0_io_coef_mainch_drc_th),
    .io_coef_mainch_drc_offset(mac_units_0_io_coef_mainch_drc_offset),
    .io_coef_mainch_drc_drcen(mac_units_0_io_coef_mainch_drc_drcen)
  );
  MacUnit mac_units_1 ( // @[dsptop.scala 88:70]
    .clock(mac_units_1_clock),
    .reset(mac_units_1_reset),
    .io_uopin_ready(mac_units_1_io_uopin_ready),
    .io_uopin_valid(mac_units_1_io_uopin_valid),
    .io_uopin_bits_vlen(mac_units_1_io_uopin_bits_vlen),
    .io_uopin_bits_select(mac_units_1_io_uopin_bits_select),
    .io_uopin_bits_drc(mac_units_1_io_uopin_bits_drc),
    .io_uopin_bits_pow(mac_units_1_io_uopin_bits_pow),
    .io_uopin_bits_loop(mac_units_1_io_uopin_bits_loop),
    .io_uopin_bits_drcgain(mac_units_1_io_uopin_bits_drcgain),
    .io_uopin_bits_drcnum(mac_units_1_io_uopin_bits_drcnum),
    .io_uopin_bits_srcreq_0_valid(mac_units_1_io_uopin_bits_srcreq_0_valid),
    .io_uopin_bits_srcreq_0_isgroup(mac_units_1_io_uopin_bits_srcreq_0_isgroup),
    .io_uopin_bits_srcreq_0_iscoef(mac_units_1_io_uopin_bits_srcreq_0_iscoef),
    .io_uopin_bits_srcreq_0_idx(mac_units_1_io_uopin_bits_srcreq_0_idx),
    .io_uopin_bits_srcreq_0_busy(mac_units_1_io_uopin_bits_srcreq_0_busy),
    .io_uopin_bits_srcreq_0_wkupidx_0(mac_units_1_io_uopin_bits_srcreq_0_wkupidx_0),
    .io_uopin_bits_srcreq_0_wkupidx_1(mac_units_1_io_uopin_bits_srcreq_0_wkupidx_1),
    .io_uopin_bits_srcreq_0_wkupidx_2(mac_units_1_io_uopin_bits_srcreq_0_wkupidx_2),
    .io_uopin_bits_srcreq_0_wkupidx_3(mac_units_1_io_uopin_bits_srcreq_0_wkupidx_3),
    .io_uopin_bits_srcreq_0_wkupidx_4(mac_units_1_io_uopin_bits_srcreq_0_wkupidx_4),
    .io_uopin_bits_srcreq_0_wkupidx_5(mac_units_1_io_uopin_bits_srcreq_0_wkupidx_5),
    .io_uopin_bits_srcreq_1_valid(mac_units_1_io_uopin_bits_srcreq_1_valid),
    .io_uopin_bits_srcreq_1_isgroup(mac_units_1_io_uopin_bits_srcreq_1_isgroup),
    .io_uopin_bits_srcreq_1_iscoef(mac_units_1_io_uopin_bits_srcreq_1_iscoef),
    .io_uopin_bits_srcreq_1_idx(mac_units_1_io_uopin_bits_srcreq_1_idx),
    .io_uopin_bits_srcreq_1_busy(mac_units_1_io_uopin_bits_srcreq_1_busy),
    .io_uopin_bits_srcreq_1_wkupidx_0(mac_units_1_io_uopin_bits_srcreq_1_wkupidx_0),
    .io_uopin_bits_srcreq_1_wkupidx_1(mac_units_1_io_uopin_bits_srcreq_1_wkupidx_1),
    .io_uopin_bits_srcreq_1_wkupidx_2(mac_units_1_io_uopin_bits_srcreq_1_wkupidx_2),
    .io_uopin_bits_srcreq_1_wkupidx_3(mac_units_1_io_uopin_bits_srcreq_1_wkupidx_3),
    .io_uopin_bits_srcreq_1_wkupidx_4(mac_units_1_io_uopin_bits_srcreq_1_wkupidx_4),
    .io_uopin_bits_srcreq_1_wkupidx_5(mac_units_1_io_uopin_bits_srcreq_1_wkupidx_5),
    .io_uopin_bits_srcreq_2_valid(mac_units_1_io_uopin_bits_srcreq_2_valid),
    .io_uopin_bits_srcreq_2_isgroup(mac_units_1_io_uopin_bits_srcreq_2_isgroup),
    .io_uopin_bits_srcreq_2_iscoef(mac_units_1_io_uopin_bits_srcreq_2_iscoef),
    .io_uopin_bits_srcreq_2_idx(mac_units_1_io_uopin_bits_srcreq_2_idx),
    .io_uopin_bits_srcreq_2_busy(mac_units_1_io_uopin_bits_srcreq_2_busy),
    .io_uopin_bits_srcreq_2_wkupidx_0(mac_units_1_io_uopin_bits_srcreq_2_wkupidx_0),
    .io_uopin_bits_srcreq_2_wkupidx_1(mac_units_1_io_uopin_bits_srcreq_2_wkupidx_1),
    .io_uopin_bits_srcreq_2_wkupidx_2(mac_units_1_io_uopin_bits_srcreq_2_wkupidx_2),
    .io_uopin_bits_srcreq_2_wkupidx_3(mac_units_1_io_uopin_bits_srcreq_2_wkupidx_3),
    .io_uopin_bits_srcreq_2_wkupidx_4(mac_units_1_io_uopin_bits_srcreq_2_wkupidx_4),
    .io_uopin_bits_srcreq_2_wkupidx_5(mac_units_1_io_uopin_bits_srcreq_2_wkupidx_5),
    .io_uopin_bits_srcreq_3_valid(mac_units_1_io_uopin_bits_srcreq_3_valid),
    .io_uopin_bits_srcreq_3_isgroup(mac_units_1_io_uopin_bits_srcreq_3_isgroup),
    .io_uopin_bits_srcreq_3_iscoef(mac_units_1_io_uopin_bits_srcreq_3_iscoef),
    .io_uopin_bits_srcreq_3_idx(mac_units_1_io_uopin_bits_srcreq_3_idx),
    .io_uopin_bits_srcreq_3_busy(mac_units_1_io_uopin_bits_srcreq_3_busy),
    .io_uopin_bits_srcreq_3_wkupidx_0(mac_units_1_io_uopin_bits_srcreq_3_wkupidx_0),
    .io_uopin_bits_srcreq_3_wkupidx_1(mac_units_1_io_uopin_bits_srcreq_3_wkupidx_1),
    .io_uopin_bits_srcreq_3_wkupidx_2(mac_units_1_io_uopin_bits_srcreq_3_wkupidx_2),
    .io_uopin_bits_srcreq_3_wkupidx_3(mac_units_1_io_uopin_bits_srcreq_3_wkupidx_3),
    .io_uopin_bits_srcreq_3_wkupidx_4(mac_units_1_io_uopin_bits_srcreq_3_wkupidx_4),
    .io_uopin_bits_srcreq_3_wkupidx_5(mac_units_1_io_uopin_bits_srcreq_3_wkupidx_5),
    .io_uopin_bits_srcreq_4_valid(mac_units_1_io_uopin_bits_srcreq_4_valid),
    .io_uopin_bits_srcreq_4_isgroup(mac_units_1_io_uopin_bits_srcreq_4_isgroup),
    .io_uopin_bits_srcreq_4_iscoef(mac_units_1_io_uopin_bits_srcreq_4_iscoef),
    .io_uopin_bits_srcreq_4_idx(mac_units_1_io_uopin_bits_srcreq_4_idx),
    .io_uopin_bits_srcreq_4_busy(mac_units_1_io_uopin_bits_srcreq_4_busy),
    .io_uopin_bits_srcreq_4_wkupidx_0(mac_units_1_io_uopin_bits_srcreq_4_wkupidx_0),
    .io_uopin_bits_srcreq_4_wkupidx_1(mac_units_1_io_uopin_bits_srcreq_4_wkupidx_1),
    .io_uopin_bits_srcreq_4_wkupidx_2(mac_units_1_io_uopin_bits_srcreq_4_wkupidx_2),
    .io_uopin_bits_srcreq_4_wkupidx_3(mac_units_1_io_uopin_bits_srcreq_4_wkupidx_3),
    .io_uopin_bits_srcreq_4_wkupidx_4(mac_units_1_io_uopin_bits_srcreq_4_wkupidx_4),
    .io_uopin_bits_srcreq_4_wkupidx_5(mac_units_1_io_uopin_bits_srcreq_4_wkupidx_5),
    .io_uopin_bits_srcreq_5_valid(mac_units_1_io_uopin_bits_srcreq_5_valid),
    .io_uopin_bits_srcreq_5_isgroup(mac_units_1_io_uopin_bits_srcreq_5_isgroup),
    .io_uopin_bits_srcreq_5_iscoef(mac_units_1_io_uopin_bits_srcreq_5_iscoef),
    .io_uopin_bits_srcreq_5_idx(mac_units_1_io_uopin_bits_srcreq_5_idx),
    .io_uopin_bits_srcreq_5_busy(mac_units_1_io_uopin_bits_srcreq_5_busy),
    .io_uopin_bits_srcreq_5_wkupidx_0(mac_units_1_io_uopin_bits_srcreq_5_wkupidx_0),
    .io_uopin_bits_srcreq_5_wkupidx_1(mac_units_1_io_uopin_bits_srcreq_5_wkupidx_1),
    .io_uopin_bits_srcreq_5_wkupidx_2(mac_units_1_io_uopin_bits_srcreq_5_wkupidx_2),
    .io_uopin_bits_srcreq_5_wkupidx_3(mac_units_1_io_uopin_bits_srcreq_5_wkupidx_3),
    .io_uopin_bits_srcreq_5_wkupidx_4(mac_units_1_io_uopin_bits_srcreq_5_wkupidx_4),
    .io_uopin_bits_srcreq_5_wkupidx_5(mac_units_1_io_uopin_bits_srcreq_5_wkupidx_5),
    .io_uopin_bits_wbvld(mac_units_1_io_uopin_bits_wbvld),
    .io_uopin_bits_wbreq(mac_units_1_io_uopin_bits_wbreq),
    .io_uopin_bits_waridx_0(mac_units_1_io_uopin_bits_waridx_0),
    .io_uopin_bits_waridx_1(mac_units_1_io_uopin_bits_waridx_1),
    .io_uopin_bits_waridx_2(mac_units_1_io_uopin_bits_waridx_2),
    .io_uopin_bits_waridx_3(mac_units_1_io_uopin_bits_waridx_3),
    .io_uopin_bits_waridx_4(mac_units_1_io_uopin_bits_waridx_4),
    .io_uopin_bits_wawidx_0(mac_units_1_io_uopin_bits_wawidx_0),
    .io_uopin_bits_wawidx_1(mac_units_1_io_uopin_bits_wawidx_1),
    .io_uopin_bits_wawidx_2(mac_units_1_io_uopin_bits_wawidx_2),
    .io_uopin_bits_wawidx_3(mac_units_1_io_uopin_bits_wawidx_3),
    .io_uopin_bits_wawidx_4(mac_units_1_io_uopin_bits_wawidx_4),
    .io_rfreq_0_req_isgroup(mac_units_1_io_rfreq_0_req_isgroup),
    .io_rfreq_0_req_iscoef(mac_units_1_io_rfreq_0_req_iscoef),
    .io_rfreq_0_req_idx(mac_units_1_io_rfreq_0_req_idx),
    .io_rfreq_0_req_gidx(mac_units_1_io_rfreq_0_req_gidx),
    .io_rfreq_0_resp(mac_units_1_io_rfreq_0_resp),
    .io_rfreq_1_req_isgroup(mac_units_1_io_rfreq_1_req_isgroup),
    .io_rfreq_1_req_iscoef(mac_units_1_io_rfreq_1_req_iscoef),
    .io_rfreq_1_req_idx(mac_units_1_io_rfreq_1_req_idx),
    .io_rfreq_1_req_gidx(mac_units_1_io_rfreq_1_req_gidx),
    .io_rfreq_1_req_sel(mac_units_1_io_rfreq_1_req_sel),
    .io_rfreq_1_resp(mac_units_1_io_rfreq_1_resp),
    .io_wbreq_wdata1(mac_units_1_io_wbreq_wdata1),
    .io_wbreq_wdata2(mac_units_1_io_wbreq_wdata2),
    .io_wbreq_vld(mac_units_1_io_wbreq_vld),
    .io_wbreq_gregidx(mac_units_1_io_wbreq_gregidx),
    .io_fwd_wkup_valid(mac_units_1_io_fwd_wkup_valid),
    .io_fwd_wkup_bits(mac_units_1_io_fwd_wkup_bits),
    .io_empty(mac_units_1_io_empty),
    .io_raw_wkup_0_valid(mac_units_1_io_raw_wkup_0_valid),
    .io_raw_wkup_0_bits(mac_units_1_io_raw_wkup_0_bits),
    .io_raw_wkup_1_valid(mac_units_1_io_raw_wkup_1_valid),
    .io_raw_wkup_1_bits(mac_units_1_io_raw_wkup_1_bits),
    .io_raw_wkup_2_valid(mac_units_1_io_raw_wkup_2_valid),
    .io_raw_wkup_2_bits(mac_units_1_io_raw_wkup_2_bits),
    .io_raw_wkup_3_valid(mac_units_1_io_raw_wkup_3_valid),
    .io_raw_wkup_3_bits(mac_units_1_io_raw_wkup_3_bits),
    .io_raw_wkup_4_valid(mac_units_1_io_raw_wkup_4_valid),
    .io_raw_wkup_4_bits(mac_units_1_io_raw_wkup_4_bits),
    .io_raw_wkup_5_valid(mac_units_1_io_raw_wkup_5_valid),
    .io_raw_wkup_5_bits(mac_units_1_io_raw_wkup_5_bits),
    .io_wbcheck_valid(mac_units_1_io_wbcheck_valid),
    .io_wbcheck_bits(mac_units_1_io_wbcheck_bits),
    .io_r_check_0_valid(mac_units_1_io_r_check_0_valid),
    .io_r_check_0_bits(mac_units_1_io_r_check_0_bits),
    .io_r_check_1_valid(mac_units_1_io_r_check_1_valid),
    .io_r_check_1_bits(mac_units_1_io_r_check_1_bits),
    .io_r_check_2_valid(mac_units_1_io_r_check_2_valid),
    .io_r_check_2_bits(mac_units_1_io_r_check_2_bits),
    .io_r_check_3_valid(mac_units_1_io_r_check_3_valid),
    .io_r_check_3_bits(mac_units_1_io_r_check_3_bits),
    .io_r_check_4_valid(mac_units_1_io_r_check_4_valid),
    .io_r_check_4_bits(mac_units_1_io_r_check_4_bits),
    .io_r_check_5_valid(mac_units_1_io_r_check_5_valid),
    .io_r_check_5_bits(mac_units_1_io_r_check_5_bits),
    .io_other_flop_0(mac_units_1_io_other_flop_0),
    .io_other_flop_1(mac_units_1_io_other_flop_1),
    .io_other_flop_2(mac_units_1_io_other_flop_2),
    .io_other_flop_3(mac_units_1_io_other_flop_3),
    .io_other_flop_4(mac_units_1_io_other_flop_4),
    .io_flop(mac_units_1_io_flop),
    .io_coef_subch_drc_th(mac_units_1_io_coef_subch_drc_th),
    .io_coef_subch_drc_offset(mac_units_1_io_coef_subch_drc_offset),
    .io_coef_subch_drc_drcen(mac_units_1_io_coef_subch_drc_drcen),
    .io_coef_mainch_ch0_autoloop(mac_units_1_io_coef_mainch_ch0_autoloop),
    .io_coef_mainch_drc_th(mac_units_1_io_coef_mainch_drc_th),
    .io_coef_mainch_drc_offset(mac_units_1_io_coef_mainch_drc_offset),
    .io_coef_mainch_drc_drcen(mac_units_1_io_coef_mainch_drc_drcen)
  );
  MacUnit mac_units_2 ( // @[dsptop.scala 88:70]
    .clock(mac_units_2_clock),
    .reset(mac_units_2_reset),
    .io_uopin_ready(mac_units_2_io_uopin_ready),
    .io_uopin_valid(mac_units_2_io_uopin_valid),
    .io_uopin_bits_vlen(mac_units_2_io_uopin_bits_vlen),
    .io_uopin_bits_select(mac_units_2_io_uopin_bits_select),
    .io_uopin_bits_drc(mac_units_2_io_uopin_bits_drc),
    .io_uopin_bits_pow(mac_units_2_io_uopin_bits_pow),
    .io_uopin_bits_loop(mac_units_2_io_uopin_bits_loop),
    .io_uopin_bits_drcgain(mac_units_2_io_uopin_bits_drcgain),
    .io_uopin_bits_drcnum(mac_units_2_io_uopin_bits_drcnum),
    .io_uopin_bits_srcreq_0_valid(mac_units_2_io_uopin_bits_srcreq_0_valid),
    .io_uopin_bits_srcreq_0_isgroup(mac_units_2_io_uopin_bits_srcreq_0_isgroup),
    .io_uopin_bits_srcreq_0_iscoef(mac_units_2_io_uopin_bits_srcreq_0_iscoef),
    .io_uopin_bits_srcreq_0_idx(mac_units_2_io_uopin_bits_srcreq_0_idx),
    .io_uopin_bits_srcreq_0_busy(mac_units_2_io_uopin_bits_srcreq_0_busy),
    .io_uopin_bits_srcreq_0_wkupidx_0(mac_units_2_io_uopin_bits_srcreq_0_wkupidx_0),
    .io_uopin_bits_srcreq_0_wkupidx_1(mac_units_2_io_uopin_bits_srcreq_0_wkupidx_1),
    .io_uopin_bits_srcreq_0_wkupidx_2(mac_units_2_io_uopin_bits_srcreq_0_wkupidx_2),
    .io_uopin_bits_srcreq_0_wkupidx_3(mac_units_2_io_uopin_bits_srcreq_0_wkupidx_3),
    .io_uopin_bits_srcreq_0_wkupidx_4(mac_units_2_io_uopin_bits_srcreq_0_wkupidx_4),
    .io_uopin_bits_srcreq_0_wkupidx_5(mac_units_2_io_uopin_bits_srcreq_0_wkupidx_5),
    .io_uopin_bits_srcreq_1_valid(mac_units_2_io_uopin_bits_srcreq_1_valid),
    .io_uopin_bits_srcreq_1_isgroup(mac_units_2_io_uopin_bits_srcreq_1_isgroup),
    .io_uopin_bits_srcreq_1_iscoef(mac_units_2_io_uopin_bits_srcreq_1_iscoef),
    .io_uopin_bits_srcreq_1_idx(mac_units_2_io_uopin_bits_srcreq_1_idx),
    .io_uopin_bits_srcreq_1_busy(mac_units_2_io_uopin_bits_srcreq_1_busy),
    .io_uopin_bits_srcreq_1_wkupidx_0(mac_units_2_io_uopin_bits_srcreq_1_wkupidx_0),
    .io_uopin_bits_srcreq_1_wkupidx_1(mac_units_2_io_uopin_bits_srcreq_1_wkupidx_1),
    .io_uopin_bits_srcreq_1_wkupidx_2(mac_units_2_io_uopin_bits_srcreq_1_wkupidx_2),
    .io_uopin_bits_srcreq_1_wkupidx_3(mac_units_2_io_uopin_bits_srcreq_1_wkupidx_3),
    .io_uopin_bits_srcreq_1_wkupidx_4(mac_units_2_io_uopin_bits_srcreq_1_wkupidx_4),
    .io_uopin_bits_srcreq_1_wkupidx_5(mac_units_2_io_uopin_bits_srcreq_1_wkupidx_5),
    .io_uopin_bits_srcreq_2_valid(mac_units_2_io_uopin_bits_srcreq_2_valid),
    .io_uopin_bits_srcreq_2_isgroup(mac_units_2_io_uopin_bits_srcreq_2_isgroup),
    .io_uopin_bits_srcreq_2_iscoef(mac_units_2_io_uopin_bits_srcreq_2_iscoef),
    .io_uopin_bits_srcreq_2_idx(mac_units_2_io_uopin_bits_srcreq_2_idx),
    .io_uopin_bits_srcreq_2_busy(mac_units_2_io_uopin_bits_srcreq_2_busy),
    .io_uopin_bits_srcreq_2_wkupidx_0(mac_units_2_io_uopin_bits_srcreq_2_wkupidx_0),
    .io_uopin_bits_srcreq_2_wkupidx_1(mac_units_2_io_uopin_bits_srcreq_2_wkupidx_1),
    .io_uopin_bits_srcreq_2_wkupidx_2(mac_units_2_io_uopin_bits_srcreq_2_wkupidx_2),
    .io_uopin_bits_srcreq_2_wkupidx_3(mac_units_2_io_uopin_bits_srcreq_2_wkupidx_3),
    .io_uopin_bits_srcreq_2_wkupidx_4(mac_units_2_io_uopin_bits_srcreq_2_wkupidx_4),
    .io_uopin_bits_srcreq_2_wkupidx_5(mac_units_2_io_uopin_bits_srcreq_2_wkupidx_5),
    .io_uopin_bits_srcreq_3_valid(mac_units_2_io_uopin_bits_srcreq_3_valid),
    .io_uopin_bits_srcreq_3_isgroup(mac_units_2_io_uopin_bits_srcreq_3_isgroup),
    .io_uopin_bits_srcreq_3_iscoef(mac_units_2_io_uopin_bits_srcreq_3_iscoef),
    .io_uopin_bits_srcreq_3_idx(mac_units_2_io_uopin_bits_srcreq_3_idx),
    .io_uopin_bits_srcreq_3_busy(mac_units_2_io_uopin_bits_srcreq_3_busy),
    .io_uopin_bits_srcreq_3_wkupidx_0(mac_units_2_io_uopin_bits_srcreq_3_wkupidx_0),
    .io_uopin_bits_srcreq_3_wkupidx_1(mac_units_2_io_uopin_bits_srcreq_3_wkupidx_1),
    .io_uopin_bits_srcreq_3_wkupidx_2(mac_units_2_io_uopin_bits_srcreq_3_wkupidx_2),
    .io_uopin_bits_srcreq_3_wkupidx_3(mac_units_2_io_uopin_bits_srcreq_3_wkupidx_3),
    .io_uopin_bits_srcreq_3_wkupidx_4(mac_units_2_io_uopin_bits_srcreq_3_wkupidx_4),
    .io_uopin_bits_srcreq_3_wkupidx_5(mac_units_2_io_uopin_bits_srcreq_3_wkupidx_5),
    .io_uopin_bits_srcreq_4_valid(mac_units_2_io_uopin_bits_srcreq_4_valid),
    .io_uopin_bits_srcreq_4_isgroup(mac_units_2_io_uopin_bits_srcreq_4_isgroup),
    .io_uopin_bits_srcreq_4_iscoef(mac_units_2_io_uopin_bits_srcreq_4_iscoef),
    .io_uopin_bits_srcreq_4_idx(mac_units_2_io_uopin_bits_srcreq_4_idx),
    .io_uopin_bits_srcreq_4_busy(mac_units_2_io_uopin_bits_srcreq_4_busy),
    .io_uopin_bits_srcreq_4_wkupidx_0(mac_units_2_io_uopin_bits_srcreq_4_wkupidx_0),
    .io_uopin_bits_srcreq_4_wkupidx_1(mac_units_2_io_uopin_bits_srcreq_4_wkupidx_1),
    .io_uopin_bits_srcreq_4_wkupidx_2(mac_units_2_io_uopin_bits_srcreq_4_wkupidx_2),
    .io_uopin_bits_srcreq_4_wkupidx_3(mac_units_2_io_uopin_bits_srcreq_4_wkupidx_3),
    .io_uopin_bits_srcreq_4_wkupidx_4(mac_units_2_io_uopin_bits_srcreq_4_wkupidx_4),
    .io_uopin_bits_srcreq_4_wkupidx_5(mac_units_2_io_uopin_bits_srcreq_4_wkupidx_5),
    .io_uopin_bits_srcreq_5_valid(mac_units_2_io_uopin_bits_srcreq_5_valid),
    .io_uopin_bits_srcreq_5_isgroup(mac_units_2_io_uopin_bits_srcreq_5_isgroup),
    .io_uopin_bits_srcreq_5_iscoef(mac_units_2_io_uopin_bits_srcreq_5_iscoef),
    .io_uopin_bits_srcreq_5_idx(mac_units_2_io_uopin_bits_srcreq_5_idx),
    .io_uopin_bits_srcreq_5_busy(mac_units_2_io_uopin_bits_srcreq_5_busy),
    .io_uopin_bits_srcreq_5_wkupidx_0(mac_units_2_io_uopin_bits_srcreq_5_wkupidx_0),
    .io_uopin_bits_srcreq_5_wkupidx_1(mac_units_2_io_uopin_bits_srcreq_5_wkupidx_1),
    .io_uopin_bits_srcreq_5_wkupidx_2(mac_units_2_io_uopin_bits_srcreq_5_wkupidx_2),
    .io_uopin_bits_srcreq_5_wkupidx_3(mac_units_2_io_uopin_bits_srcreq_5_wkupidx_3),
    .io_uopin_bits_srcreq_5_wkupidx_4(mac_units_2_io_uopin_bits_srcreq_5_wkupidx_4),
    .io_uopin_bits_srcreq_5_wkupidx_5(mac_units_2_io_uopin_bits_srcreq_5_wkupidx_5),
    .io_uopin_bits_wbvld(mac_units_2_io_uopin_bits_wbvld),
    .io_uopin_bits_wbreq(mac_units_2_io_uopin_bits_wbreq),
    .io_uopin_bits_waridx_0(mac_units_2_io_uopin_bits_waridx_0),
    .io_uopin_bits_waridx_1(mac_units_2_io_uopin_bits_waridx_1),
    .io_uopin_bits_waridx_2(mac_units_2_io_uopin_bits_waridx_2),
    .io_uopin_bits_waridx_3(mac_units_2_io_uopin_bits_waridx_3),
    .io_uopin_bits_waridx_4(mac_units_2_io_uopin_bits_waridx_4),
    .io_uopin_bits_wawidx_0(mac_units_2_io_uopin_bits_wawidx_0),
    .io_uopin_bits_wawidx_1(mac_units_2_io_uopin_bits_wawidx_1),
    .io_uopin_bits_wawidx_2(mac_units_2_io_uopin_bits_wawidx_2),
    .io_uopin_bits_wawidx_3(mac_units_2_io_uopin_bits_wawidx_3),
    .io_uopin_bits_wawidx_4(mac_units_2_io_uopin_bits_wawidx_4),
    .io_rfreq_0_req_isgroup(mac_units_2_io_rfreq_0_req_isgroup),
    .io_rfreq_0_req_iscoef(mac_units_2_io_rfreq_0_req_iscoef),
    .io_rfreq_0_req_idx(mac_units_2_io_rfreq_0_req_idx),
    .io_rfreq_0_req_gidx(mac_units_2_io_rfreq_0_req_gidx),
    .io_rfreq_0_resp(mac_units_2_io_rfreq_0_resp),
    .io_rfreq_1_req_isgroup(mac_units_2_io_rfreq_1_req_isgroup),
    .io_rfreq_1_req_iscoef(mac_units_2_io_rfreq_1_req_iscoef),
    .io_rfreq_1_req_idx(mac_units_2_io_rfreq_1_req_idx),
    .io_rfreq_1_req_gidx(mac_units_2_io_rfreq_1_req_gidx),
    .io_rfreq_1_req_sel(mac_units_2_io_rfreq_1_req_sel),
    .io_rfreq_1_resp(mac_units_2_io_rfreq_1_resp),
    .io_wbreq_wdata1(mac_units_2_io_wbreq_wdata1),
    .io_wbreq_wdata2(mac_units_2_io_wbreq_wdata2),
    .io_wbreq_vld(mac_units_2_io_wbreq_vld),
    .io_wbreq_gregidx(mac_units_2_io_wbreq_gregidx),
    .io_fwd_wkup_valid(mac_units_2_io_fwd_wkup_valid),
    .io_fwd_wkup_bits(mac_units_2_io_fwd_wkup_bits),
    .io_empty(mac_units_2_io_empty),
    .io_raw_wkup_0_valid(mac_units_2_io_raw_wkup_0_valid),
    .io_raw_wkup_0_bits(mac_units_2_io_raw_wkup_0_bits),
    .io_raw_wkup_1_valid(mac_units_2_io_raw_wkup_1_valid),
    .io_raw_wkup_1_bits(mac_units_2_io_raw_wkup_1_bits),
    .io_raw_wkup_2_valid(mac_units_2_io_raw_wkup_2_valid),
    .io_raw_wkup_2_bits(mac_units_2_io_raw_wkup_2_bits),
    .io_raw_wkup_3_valid(mac_units_2_io_raw_wkup_3_valid),
    .io_raw_wkup_3_bits(mac_units_2_io_raw_wkup_3_bits),
    .io_raw_wkup_4_valid(mac_units_2_io_raw_wkup_4_valid),
    .io_raw_wkup_4_bits(mac_units_2_io_raw_wkup_4_bits),
    .io_raw_wkup_5_valid(mac_units_2_io_raw_wkup_5_valid),
    .io_raw_wkup_5_bits(mac_units_2_io_raw_wkup_5_bits),
    .io_wbcheck_valid(mac_units_2_io_wbcheck_valid),
    .io_wbcheck_bits(mac_units_2_io_wbcheck_bits),
    .io_r_check_0_valid(mac_units_2_io_r_check_0_valid),
    .io_r_check_0_bits(mac_units_2_io_r_check_0_bits),
    .io_r_check_1_valid(mac_units_2_io_r_check_1_valid),
    .io_r_check_1_bits(mac_units_2_io_r_check_1_bits),
    .io_r_check_2_valid(mac_units_2_io_r_check_2_valid),
    .io_r_check_2_bits(mac_units_2_io_r_check_2_bits),
    .io_r_check_3_valid(mac_units_2_io_r_check_3_valid),
    .io_r_check_3_bits(mac_units_2_io_r_check_3_bits),
    .io_r_check_4_valid(mac_units_2_io_r_check_4_valid),
    .io_r_check_4_bits(mac_units_2_io_r_check_4_bits),
    .io_r_check_5_valid(mac_units_2_io_r_check_5_valid),
    .io_r_check_5_bits(mac_units_2_io_r_check_5_bits),
    .io_other_flop_0(mac_units_2_io_other_flop_0),
    .io_other_flop_1(mac_units_2_io_other_flop_1),
    .io_other_flop_2(mac_units_2_io_other_flop_2),
    .io_other_flop_3(mac_units_2_io_other_flop_3),
    .io_other_flop_4(mac_units_2_io_other_flop_4),
    .io_flop(mac_units_2_io_flop),
    .io_coef_subch_drc_th(mac_units_2_io_coef_subch_drc_th),
    .io_coef_subch_drc_offset(mac_units_2_io_coef_subch_drc_offset),
    .io_coef_subch_drc_drcen(mac_units_2_io_coef_subch_drc_drcen),
    .io_coef_mainch_ch0_autoloop(mac_units_2_io_coef_mainch_ch0_autoloop),
    .io_coef_mainch_drc_th(mac_units_2_io_coef_mainch_drc_th),
    .io_coef_mainch_drc_offset(mac_units_2_io_coef_mainch_drc_offset),
    .io_coef_mainch_drc_drcen(mac_units_2_io_coef_mainch_drc_drcen)
  );
  MacUnit mac_units_3 ( // @[dsptop.scala 88:70]
    .clock(mac_units_3_clock),
    .reset(mac_units_3_reset),
    .io_uopin_ready(mac_units_3_io_uopin_ready),
    .io_uopin_valid(mac_units_3_io_uopin_valid),
    .io_uopin_bits_vlen(mac_units_3_io_uopin_bits_vlen),
    .io_uopin_bits_select(mac_units_3_io_uopin_bits_select),
    .io_uopin_bits_drc(mac_units_3_io_uopin_bits_drc),
    .io_uopin_bits_pow(mac_units_3_io_uopin_bits_pow),
    .io_uopin_bits_loop(mac_units_3_io_uopin_bits_loop),
    .io_uopin_bits_drcgain(mac_units_3_io_uopin_bits_drcgain),
    .io_uopin_bits_drcnum(mac_units_3_io_uopin_bits_drcnum),
    .io_uopin_bits_srcreq_0_valid(mac_units_3_io_uopin_bits_srcreq_0_valid),
    .io_uopin_bits_srcreq_0_isgroup(mac_units_3_io_uopin_bits_srcreq_0_isgroup),
    .io_uopin_bits_srcreq_0_iscoef(mac_units_3_io_uopin_bits_srcreq_0_iscoef),
    .io_uopin_bits_srcreq_0_idx(mac_units_3_io_uopin_bits_srcreq_0_idx),
    .io_uopin_bits_srcreq_0_busy(mac_units_3_io_uopin_bits_srcreq_0_busy),
    .io_uopin_bits_srcreq_0_wkupidx_0(mac_units_3_io_uopin_bits_srcreq_0_wkupidx_0),
    .io_uopin_bits_srcreq_0_wkupidx_1(mac_units_3_io_uopin_bits_srcreq_0_wkupidx_1),
    .io_uopin_bits_srcreq_0_wkupidx_2(mac_units_3_io_uopin_bits_srcreq_0_wkupidx_2),
    .io_uopin_bits_srcreq_0_wkupidx_3(mac_units_3_io_uopin_bits_srcreq_0_wkupidx_3),
    .io_uopin_bits_srcreq_0_wkupidx_4(mac_units_3_io_uopin_bits_srcreq_0_wkupidx_4),
    .io_uopin_bits_srcreq_0_wkupidx_5(mac_units_3_io_uopin_bits_srcreq_0_wkupidx_5),
    .io_uopin_bits_srcreq_1_valid(mac_units_3_io_uopin_bits_srcreq_1_valid),
    .io_uopin_bits_srcreq_1_isgroup(mac_units_3_io_uopin_bits_srcreq_1_isgroup),
    .io_uopin_bits_srcreq_1_iscoef(mac_units_3_io_uopin_bits_srcreq_1_iscoef),
    .io_uopin_bits_srcreq_1_idx(mac_units_3_io_uopin_bits_srcreq_1_idx),
    .io_uopin_bits_srcreq_1_busy(mac_units_3_io_uopin_bits_srcreq_1_busy),
    .io_uopin_bits_srcreq_1_wkupidx_0(mac_units_3_io_uopin_bits_srcreq_1_wkupidx_0),
    .io_uopin_bits_srcreq_1_wkupidx_1(mac_units_3_io_uopin_bits_srcreq_1_wkupidx_1),
    .io_uopin_bits_srcreq_1_wkupidx_2(mac_units_3_io_uopin_bits_srcreq_1_wkupidx_2),
    .io_uopin_bits_srcreq_1_wkupidx_3(mac_units_3_io_uopin_bits_srcreq_1_wkupidx_3),
    .io_uopin_bits_srcreq_1_wkupidx_4(mac_units_3_io_uopin_bits_srcreq_1_wkupidx_4),
    .io_uopin_bits_srcreq_1_wkupidx_5(mac_units_3_io_uopin_bits_srcreq_1_wkupidx_5),
    .io_uopin_bits_srcreq_2_valid(mac_units_3_io_uopin_bits_srcreq_2_valid),
    .io_uopin_bits_srcreq_2_isgroup(mac_units_3_io_uopin_bits_srcreq_2_isgroup),
    .io_uopin_bits_srcreq_2_iscoef(mac_units_3_io_uopin_bits_srcreq_2_iscoef),
    .io_uopin_bits_srcreq_2_idx(mac_units_3_io_uopin_bits_srcreq_2_idx),
    .io_uopin_bits_srcreq_2_busy(mac_units_3_io_uopin_bits_srcreq_2_busy),
    .io_uopin_bits_srcreq_2_wkupidx_0(mac_units_3_io_uopin_bits_srcreq_2_wkupidx_0),
    .io_uopin_bits_srcreq_2_wkupidx_1(mac_units_3_io_uopin_bits_srcreq_2_wkupidx_1),
    .io_uopin_bits_srcreq_2_wkupidx_2(mac_units_3_io_uopin_bits_srcreq_2_wkupidx_2),
    .io_uopin_bits_srcreq_2_wkupidx_3(mac_units_3_io_uopin_bits_srcreq_2_wkupidx_3),
    .io_uopin_bits_srcreq_2_wkupidx_4(mac_units_3_io_uopin_bits_srcreq_2_wkupidx_4),
    .io_uopin_bits_srcreq_2_wkupidx_5(mac_units_3_io_uopin_bits_srcreq_2_wkupidx_5),
    .io_uopin_bits_srcreq_3_valid(mac_units_3_io_uopin_bits_srcreq_3_valid),
    .io_uopin_bits_srcreq_3_isgroup(mac_units_3_io_uopin_bits_srcreq_3_isgroup),
    .io_uopin_bits_srcreq_3_iscoef(mac_units_3_io_uopin_bits_srcreq_3_iscoef),
    .io_uopin_bits_srcreq_3_idx(mac_units_3_io_uopin_bits_srcreq_3_idx),
    .io_uopin_bits_srcreq_3_busy(mac_units_3_io_uopin_bits_srcreq_3_busy),
    .io_uopin_bits_srcreq_3_wkupidx_0(mac_units_3_io_uopin_bits_srcreq_3_wkupidx_0),
    .io_uopin_bits_srcreq_3_wkupidx_1(mac_units_3_io_uopin_bits_srcreq_3_wkupidx_1),
    .io_uopin_bits_srcreq_3_wkupidx_2(mac_units_3_io_uopin_bits_srcreq_3_wkupidx_2),
    .io_uopin_bits_srcreq_3_wkupidx_3(mac_units_3_io_uopin_bits_srcreq_3_wkupidx_3),
    .io_uopin_bits_srcreq_3_wkupidx_4(mac_units_3_io_uopin_bits_srcreq_3_wkupidx_4),
    .io_uopin_bits_srcreq_3_wkupidx_5(mac_units_3_io_uopin_bits_srcreq_3_wkupidx_5),
    .io_uopin_bits_srcreq_4_valid(mac_units_3_io_uopin_bits_srcreq_4_valid),
    .io_uopin_bits_srcreq_4_isgroup(mac_units_3_io_uopin_bits_srcreq_4_isgroup),
    .io_uopin_bits_srcreq_4_iscoef(mac_units_3_io_uopin_bits_srcreq_4_iscoef),
    .io_uopin_bits_srcreq_4_idx(mac_units_3_io_uopin_bits_srcreq_4_idx),
    .io_uopin_bits_srcreq_4_busy(mac_units_3_io_uopin_bits_srcreq_4_busy),
    .io_uopin_bits_srcreq_4_wkupidx_0(mac_units_3_io_uopin_bits_srcreq_4_wkupidx_0),
    .io_uopin_bits_srcreq_4_wkupidx_1(mac_units_3_io_uopin_bits_srcreq_4_wkupidx_1),
    .io_uopin_bits_srcreq_4_wkupidx_2(mac_units_3_io_uopin_bits_srcreq_4_wkupidx_2),
    .io_uopin_bits_srcreq_4_wkupidx_3(mac_units_3_io_uopin_bits_srcreq_4_wkupidx_3),
    .io_uopin_bits_srcreq_4_wkupidx_4(mac_units_3_io_uopin_bits_srcreq_4_wkupidx_4),
    .io_uopin_bits_srcreq_4_wkupidx_5(mac_units_3_io_uopin_bits_srcreq_4_wkupidx_5),
    .io_uopin_bits_srcreq_5_valid(mac_units_3_io_uopin_bits_srcreq_5_valid),
    .io_uopin_bits_srcreq_5_isgroup(mac_units_3_io_uopin_bits_srcreq_5_isgroup),
    .io_uopin_bits_srcreq_5_iscoef(mac_units_3_io_uopin_bits_srcreq_5_iscoef),
    .io_uopin_bits_srcreq_5_idx(mac_units_3_io_uopin_bits_srcreq_5_idx),
    .io_uopin_bits_srcreq_5_busy(mac_units_3_io_uopin_bits_srcreq_5_busy),
    .io_uopin_bits_srcreq_5_wkupidx_0(mac_units_3_io_uopin_bits_srcreq_5_wkupidx_0),
    .io_uopin_bits_srcreq_5_wkupidx_1(mac_units_3_io_uopin_bits_srcreq_5_wkupidx_1),
    .io_uopin_bits_srcreq_5_wkupidx_2(mac_units_3_io_uopin_bits_srcreq_5_wkupidx_2),
    .io_uopin_bits_srcreq_5_wkupidx_3(mac_units_3_io_uopin_bits_srcreq_5_wkupidx_3),
    .io_uopin_bits_srcreq_5_wkupidx_4(mac_units_3_io_uopin_bits_srcreq_5_wkupidx_4),
    .io_uopin_bits_srcreq_5_wkupidx_5(mac_units_3_io_uopin_bits_srcreq_5_wkupidx_5),
    .io_uopin_bits_wbvld(mac_units_3_io_uopin_bits_wbvld),
    .io_uopin_bits_wbreq(mac_units_3_io_uopin_bits_wbreq),
    .io_uopin_bits_waridx_0(mac_units_3_io_uopin_bits_waridx_0),
    .io_uopin_bits_waridx_1(mac_units_3_io_uopin_bits_waridx_1),
    .io_uopin_bits_waridx_2(mac_units_3_io_uopin_bits_waridx_2),
    .io_uopin_bits_waridx_3(mac_units_3_io_uopin_bits_waridx_3),
    .io_uopin_bits_waridx_4(mac_units_3_io_uopin_bits_waridx_4),
    .io_uopin_bits_wawidx_0(mac_units_3_io_uopin_bits_wawidx_0),
    .io_uopin_bits_wawidx_1(mac_units_3_io_uopin_bits_wawidx_1),
    .io_uopin_bits_wawidx_2(mac_units_3_io_uopin_bits_wawidx_2),
    .io_uopin_bits_wawidx_3(mac_units_3_io_uopin_bits_wawidx_3),
    .io_uopin_bits_wawidx_4(mac_units_3_io_uopin_bits_wawidx_4),
    .io_rfreq_0_req_isgroup(mac_units_3_io_rfreq_0_req_isgroup),
    .io_rfreq_0_req_iscoef(mac_units_3_io_rfreq_0_req_iscoef),
    .io_rfreq_0_req_idx(mac_units_3_io_rfreq_0_req_idx),
    .io_rfreq_0_req_gidx(mac_units_3_io_rfreq_0_req_gidx),
    .io_rfreq_0_resp(mac_units_3_io_rfreq_0_resp),
    .io_rfreq_1_req_isgroup(mac_units_3_io_rfreq_1_req_isgroup),
    .io_rfreq_1_req_iscoef(mac_units_3_io_rfreq_1_req_iscoef),
    .io_rfreq_1_req_idx(mac_units_3_io_rfreq_1_req_idx),
    .io_rfreq_1_req_gidx(mac_units_3_io_rfreq_1_req_gidx),
    .io_rfreq_1_req_sel(mac_units_3_io_rfreq_1_req_sel),
    .io_rfreq_1_resp(mac_units_3_io_rfreq_1_resp),
    .io_wbreq_wdata1(mac_units_3_io_wbreq_wdata1),
    .io_wbreq_wdata2(mac_units_3_io_wbreq_wdata2),
    .io_wbreq_vld(mac_units_3_io_wbreq_vld),
    .io_wbreq_gregidx(mac_units_3_io_wbreq_gregidx),
    .io_fwd_wkup_valid(mac_units_3_io_fwd_wkup_valid),
    .io_fwd_wkup_bits(mac_units_3_io_fwd_wkup_bits),
    .io_empty(mac_units_3_io_empty),
    .io_raw_wkup_0_valid(mac_units_3_io_raw_wkup_0_valid),
    .io_raw_wkup_0_bits(mac_units_3_io_raw_wkup_0_bits),
    .io_raw_wkup_1_valid(mac_units_3_io_raw_wkup_1_valid),
    .io_raw_wkup_1_bits(mac_units_3_io_raw_wkup_1_bits),
    .io_raw_wkup_2_valid(mac_units_3_io_raw_wkup_2_valid),
    .io_raw_wkup_2_bits(mac_units_3_io_raw_wkup_2_bits),
    .io_raw_wkup_3_valid(mac_units_3_io_raw_wkup_3_valid),
    .io_raw_wkup_3_bits(mac_units_3_io_raw_wkup_3_bits),
    .io_raw_wkup_4_valid(mac_units_3_io_raw_wkup_4_valid),
    .io_raw_wkup_4_bits(mac_units_3_io_raw_wkup_4_bits),
    .io_raw_wkup_5_valid(mac_units_3_io_raw_wkup_5_valid),
    .io_raw_wkup_5_bits(mac_units_3_io_raw_wkup_5_bits),
    .io_wbcheck_valid(mac_units_3_io_wbcheck_valid),
    .io_wbcheck_bits(mac_units_3_io_wbcheck_bits),
    .io_r_check_0_valid(mac_units_3_io_r_check_0_valid),
    .io_r_check_0_bits(mac_units_3_io_r_check_0_bits),
    .io_r_check_1_valid(mac_units_3_io_r_check_1_valid),
    .io_r_check_1_bits(mac_units_3_io_r_check_1_bits),
    .io_r_check_2_valid(mac_units_3_io_r_check_2_valid),
    .io_r_check_2_bits(mac_units_3_io_r_check_2_bits),
    .io_r_check_3_valid(mac_units_3_io_r_check_3_valid),
    .io_r_check_3_bits(mac_units_3_io_r_check_3_bits),
    .io_r_check_4_valid(mac_units_3_io_r_check_4_valid),
    .io_r_check_4_bits(mac_units_3_io_r_check_4_bits),
    .io_r_check_5_valid(mac_units_3_io_r_check_5_valid),
    .io_r_check_5_bits(mac_units_3_io_r_check_5_bits),
    .io_other_flop_0(mac_units_3_io_other_flop_0),
    .io_other_flop_1(mac_units_3_io_other_flop_1),
    .io_other_flop_2(mac_units_3_io_other_flop_2),
    .io_other_flop_3(mac_units_3_io_other_flop_3),
    .io_other_flop_4(mac_units_3_io_other_flop_4),
    .io_flop(mac_units_3_io_flop),
    .io_coef_subch_drc_th(mac_units_3_io_coef_subch_drc_th),
    .io_coef_subch_drc_offset(mac_units_3_io_coef_subch_drc_offset),
    .io_coef_subch_drc_drcen(mac_units_3_io_coef_subch_drc_drcen),
    .io_coef_mainch_ch0_autoloop(mac_units_3_io_coef_mainch_ch0_autoloop),
    .io_coef_mainch_drc_th(mac_units_3_io_coef_mainch_drc_th),
    .io_coef_mainch_drc_offset(mac_units_3_io_coef_mainch_drc_offset),
    .io_coef_mainch_drc_drcen(mac_units_3_io_coef_mainch_drc_drcen)
  );
  MacUnit mac_units_4 ( // @[dsptop.scala 88:70]
    .clock(mac_units_4_clock),
    .reset(mac_units_4_reset),
    .io_uopin_ready(mac_units_4_io_uopin_ready),
    .io_uopin_valid(mac_units_4_io_uopin_valid),
    .io_uopin_bits_vlen(mac_units_4_io_uopin_bits_vlen),
    .io_uopin_bits_select(mac_units_4_io_uopin_bits_select),
    .io_uopin_bits_drc(mac_units_4_io_uopin_bits_drc),
    .io_uopin_bits_pow(mac_units_4_io_uopin_bits_pow),
    .io_uopin_bits_loop(mac_units_4_io_uopin_bits_loop),
    .io_uopin_bits_drcgain(mac_units_4_io_uopin_bits_drcgain),
    .io_uopin_bits_drcnum(mac_units_4_io_uopin_bits_drcnum),
    .io_uopin_bits_srcreq_0_valid(mac_units_4_io_uopin_bits_srcreq_0_valid),
    .io_uopin_bits_srcreq_0_isgroup(mac_units_4_io_uopin_bits_srcreq_0_isgroup),
    .io_uopin_bits_srcreq_0_iscoef(mac_units_4_io_uopin_bits_srcreq_0_iscoef),
    .io_uopin_bits_srcreq_0_idx(mac_units_4_io_uopin_bits_srcreq_0_idx),
    .io_uopin_bits_srcreq_0_busy(mac_units_4_io_uopin_bits_srcreq_0_busy),
    .io_uopin_bits_srcreq_0_wkupidx_0(mac_units_4_io_uopin_bits_srcreq_0_wkupidx_0),
    .io_uopin_bits_srcreq_0_wkupidx_1(mac_units_4_io_uopin_bits_srcreq_0_wkupidx_1),
    .io_uopin_bits_srcreq_0_wkupidx_2(mac_units_4_io_uopin_bits_srcreq_0_wkupidx_2),
    .io_uopin_bits_srcreq_0_wkupidx_3(mac_units_4_io_uopin_bits_srcreq_0_wkupidx_3),
    .io_uopin_bits_srcreq_0_wkupidx_4(mac_units_4_io_uopin_bits_srcreq_0_wkupidx_4),
    .io_uopin_bits_srcreq_0_wkupidx_5(mac_units_4_io_uopin_bits_srcreq_0_wkupidx_5),
    .io_uopin_bits_srcreq_1_valid(mac_units_4_io_uopin_bits_srcreq_1_valid),
    .io_uopin_bits_srcreq_1_isgroup(mac_units_4_io_uopin_bits_srcreq_1_isgroup),
    .io_uopin_bits_srcreq_1_iscoef(mac_units_4_io_uopin_bits_srcreq_1_iscoef),
    .io_uopin_bits_srcreq_1_idx(mac_units_4_io_uopin_bits_srcreq_1_idx),
    .io_uopin_bits_srcreq_1_busy(mac_units_4_io_uopin_bits_srcreq_1_busy),
    .io_uopin_bits_srcreq_1_wkupidx_0(mac_units_4_io_uopin_bits_srcreq_1_wkupidx_0),
    .io_uopin_bits_srcreq_1_wkupidx_1(mac_units_4_io_uopin_bits_srcreq_1_wkupidx_1),
    .io_uopin_bits_srcreq_1_wkupidx_2(mac_units_4_io_uopin_bits_srcreq_1_wkupidx_2),
    .io_uopin_bits_srcreq_1_wkupidx_3(mac_units_4_io_uopin_bits_srcreq_1_wkupidx_3),
    .io_uopin_bits_srcreq_1_wkupidx_4(mac_units_4_io_uopin_bits_srcreq_1_wkupidx_4),
    .io_uopin_bits_srcreq_1_wkupidx_5(mac_units_4_io_uopin_bits_srcreq_1_wkupidx_5),
    .io_uopin_bits_srcreq_2_valid(mac_units_4_io_uopin_bits_srcreq_2_valid),
    .io_uopin_bits_srcreq_2_isgroup(mac_units_4_io_uopin_bits_srcreq_2_isgroup),
    .io_uopin_bits_srcreq_2_iscoef(mac_units_4_io_uopin_bits_srcreq_2_iscoef),
    .io_uopin_bits_srcreq_2_idx(mac_units_4_io_uopin_bits_srcreq_2_idx),
    .io_uopin_bits_srcreq_2_busy(mac_units_4_io_uopin_bits_srcreq_2_busy),
    .io_uopin_bits_srcreq_2_wkupidx_0(mac_units_4_io_uopin_bits_srcreq_2_wkupidx_0),
    .io_uopin_bits_srcreq_2_wkupidx_1(mac_units_4_io_uopin_bits_srcreq_2_wkupidx_1),
    .io_uopin_bits_srcreq_2_wkupidx_2(mac_units_4_io_uopin_bits_srcreq_2_wkupidx_2),
    .io_uopin_bits_srcreq_2_wkupidx_3(mac_units_4_io_uopin_bits_srcreq_2_wkupidx_3),
    .io_uopin_bits_srcreq_2_wkupidx_4(mac_units_4_io_uopin_bits_srcreq_2_wkupidx_4),
    .io_uopin_bits_srcreq_2_wkupidx_5(mac_units_4_io_uopin_bits_srcreq_2_wkupidx_5),
    .io_uopin_bits_srcreq_3_valid(mac_units_4_io_uopin_bits_srcreq_3_valid),
    .io_uopin_bits_srcreq_3_isgroup(mac_units_4_io_uopin_bits_srcreq_3_isgroup),
    .io_uopin_bits_srcreq_3_iscoef(mac_units_4_io_uopin_bits_srcreq_3_iscoef),
    .io_uopin_bits_srcreq_3_idx(mac_units_4_io_uopin_bits_srcreq_3_idx),
    .io_uopin_bits_srcreq_3_busy(mac_units_4_io_uopin_bits_srcreq_3_busy),
    .io_uopin_bits_srcreq_3_wkupidx_0(mac_units_4_io_uopin_bits_srcreq_3_wkupidx_0),
    .io_uopin_bits_srcreq_3_wkupidx_1(mac_units_4_io_uopin_bits_srcreq_3_wkupidx_1),
    .io_uopin_bits_srcreq_3_wkupidx_2(mac_units_4_io_uopin_bits_srcreq_3_wkupidx_2),
    .io_uopin_bits_srcreq_3_wkupidx_3(mac_units_4_io_uopin_bits_srcreq_3_wkupidx_3),
    .io_uopin_bits_srcreq_3_wkupidx_4(mac_units_4_io_uopin_bits_srcreq_3_wkupidx_4),
    .io_uopin_bits_srcreq_3_wkupidx_5(mac_units_4_io_uopin_bits_srcreq_3_wkupidx_5),
    .io_uopin_bits_srcreq_4_valid(mac_units_4_io_uopin_bits_srcreq_4_valid),
    .io_uopin_bits_srcreq_4_isgroup(mac_units_4_io_uopin_bits_srcreq_4_isgroup),
    .io_uopin_bits_srcreq_4_iscoef(mac_units_4_io_uopin_bits_srcreq_4_iscoef),
    .io_uopin_bits_srcreq_4_idx(mac_units_4_io_uopin_bits_srcreq_4_idx),
    .io_uopin_bits_srcreq_4_busy(mac_units_4_io_uopin_bits_srcreq_4_busy),
    .io_uopin_bits_srcreq_4_wkupidx_0(mac_units_4_io_uopin_bits_srcreq_4_wkupidx_0),
    .io_uopin_bits_srcreq_4_wkupidx_1(mac_units_4_io_uopin_bits_srcreq_4_wkupidx_1),
    .io_uopin_bits_srcreq_4_wkupidx_2(mac_units_4_io_uopin_bits_srcreq_4_wkupidx_2),
    .io_uopin_bits_srcreq_4_wkupidx_3(mac_units_4_io_uopin_bits_srcreq_4_wkupidx_3),
    .io_uopin_bits_srcreq_4_wkupidx_4(mac_units_4_io_uopin_bits_srcreq_4_wkupidx_4),
    .io_uopin_bits_srcreq_4_wkupidx_5(mac_units_4_io_uopin_bits_srcreq_4_wkupidx_5),
    .io_uopin_bits_srcreq_5_valid(mac_units_4_io_uopin_bits_srcreq_5_valid),
    .io_uopin_bits_srcreq_5_isgroup(mac_units_4_io_uopin_bits_srcreq_5_isgroup),
    .io_uopin_bits_srcreq_5_iscoef(mac_units_4_io_uopin_bits_srcreq_5_iscoef),
    .io_uopin_bits_srcreq_5_idx(mac_units_4_io_uopin_bits_srcreq_5_idx),
    .io_uopin_bits_srcreq_5_busy(mac_units_4_io_uopin_bits_srcreq_5_busy),
    .io_uopin_bits_srcreq_5_wkupidx_0(mac_units_4_io_uopin_bits_srcreq_5_wkupidx_0),
    .io_uopin_bits_srcreq_5_wkupidx_1(mac_units_4_io_uopin_bits_srcreq_5_wkupidx_1),
    .io_uopin_bits_srcreq_5_wkupidx_2(mac_units_4_io_uopin_bits_srcreq_5_wkupidx_2),
    .io_uopin_bits_srcreq_5_wkupidx_3(mac_units_4_io_uopin_bits_srcreq_5_wkupidx_3),
    .io_uopin_bits_srcreq_5_wkupidx_4(mac_units_4_io_uopin_bits_srcreq_5_wkupidx_4),
    .io_uopin_bits_srcreq_5_wkupidx_5(mac_units_4_io_uopin_bits_srcreq_5_wkupidx_5),
    .io_uopin_bits_wbvld(mac_units_4_io_uopin_bits_wbvld),
    .io_uopin_bits_wbreq(mac_units_4_io_uopin_bits_wbreq),
    .io_uopin_bits_waridx_0(mac_units_4_io_uopin_bits_waridx_0),
    .io_uopin_bits_waridx_1(mac_units_4_io_uopin_bits_waridx_1),
    .io_uopin_bits_waridx_2(mac_units_4_io_uopin_bits_waridx_2),
    .io_uopin_bits_waridx_3(mac_units_4_io_uopin_bits_waridx_3),
    .io_uopin_bits_waridx_4(mac_units_4_io_uopin_bits_waridx_4),
    .io_uopin_bits_wawidx_0(mac_units_4_io_uopin_bits_wawidx_0),
    .io_uopin_bits_wawidx_1(mac_units_4_io_uopin_bits_wawidx_1),
    .io_uopin_bits_wawidx_2(mac_units_4_io_uopin_bits_wawidx_2),
    .io_uopin_bits_wawidx_3(mac_units_4_io_uopin_bits_wawidx_3),
    .io_uopin_bits_wawidx_4(mac_units_4_io_uopin_bits_wawidx_4),
    .io_rfreq_0_req_isgroup(mac_units_4_io_rfreq_0_req_isgroup),
    .io_rfreq_0_req_iscoef(mac_units_4_io_rfreq_0_req_iscoef),
    .io_rfreq_0_req_idx(mac_units_4_io_rfreq_0_req_idx),
    .io_rfreq_0_req_gidx(mac_units_4_io_rfreq_0_req_gidx),
    .io_rfreq_0_resp(mac_units_4_io_rfreq_0_resp),
    .io_rfreq_1_req_isgroup(mac_units_4_io_rfreq_1_req_isgroup),
    .io_rfreq_1_req_iscoef(mac_units_4_io_rfreq_1_req_iscoef),
    .io_rfreq_1_req_idx(mac_units_4_io_rfreq_1_req_idx),
    .io_rfreq_1_req_gidx(mac_units_4_io_rfreq_1_req_gidx),
    .io_rfreq_1_req_sel(mac_units_4_io_rfreq_1_req_sel),
    .io_rfreq_1_resp(mac_units_4_io_rfreq_1_resp),
    .io_wbreq_wdata1(mac_units_4_io_wbreq_wdata1),
    .io_wbreq_wdata2(mac_units_4_io_wbreq_wdata2),
    .io_wbreq_vld(mac_units_4_io_wbreq_vld),
    .io_wbreq_gregidx(mac_units_4_io_wbreq_gregidx),
    .io_fwd_wkup_valid(mac_units_4_io_fwd_wkup_valid),
    .io_fwd_wkup_bits(mac_units_4_io_fwd_wkup_bits),
    .io_empty(mac_units_4_io_empty),
    .io_raw_wkup_0_valid(mac_units_4_io_raw_wkup_0_valid),
    .io_raw_wkup_0_bits(mac_units_4_io_raw_wkup_0_bits),
    .io_raw_wkup_1_valid(mac_units_4_io_raw_wkup_1_valid),
    .io_raw_wkup_1_bits(mac_units_4_io_raw_wkup_1_bits),
    .io_raw_wkup_2_valid(mac_units_4_io_raw_wkup_2_valid),
    .io_raw_wkup_2_bits(mac_units_4_io_raw_wkup_2_bits),
    .io_raw_wkup_3_valid(mac_units_4_io_raw_wkup_3_valid),
    .io_raw_wkup_3_bits(mac_units_4_io_raw_wkup_3_bits),
    .io_raw_wkup_4_valid(mac_units_4_io_raw_wkup_4_valid),
    .io_raw_wkup_4_bits(mac_units_4_io_raw_wkup_4_bits),
    .io_raw_wkup_5_valid(mac_units_4_io_raw_wkup_5_valid),
    .io_raw_wkup_5_bits(mac_units_4_io_raw_wkup_5_bits),
    .io_wbcheck_valid(mac_units_4_io_wbcheck_valid),
    .io_wbcheck_bits(mac_units_4_io_wbcheck_bits),
    .io_r_check_0_valid(mac_units_4_io_r_check_0_valid),
    .io_r_check_0_bits(mac_units_4_io_r_check_0_bits),
    .io_r_check_1_valid(mac_units_4_io_r_check_1_valid),
    .io_r_check_1_bits(mac_units_4_io_r_check_1_bits),
    .io_r_check_2_valid(mac_units_4_io_r_check_2_valid),
    .io_r_check_2_bits(mac_units_4_io_r_check_2_bits),
    .io_r_check_3_valid(mac_units_4_io_r_check_3_valid),
    .io_r_check_3_bits(mac_units_4_io_r_check_3_bits),
    .io_r_check_4_valid(mac_units_4_io_r_check_4_valid),
    .io_r_check_4_bits(mac_units_4_io_r_check_4_bits),
    .io_r_check_5_valid(mac_units_4_io_r_check_5_valid),
    .io_r_check_5_bits(mac_units_4_io_r_check_5_bits),
    .io_other_flop_0(mac_units_4_io_other_flop_0),
    .io_other_flop_1(mac_units_4_io_other_flop_1),
    .io_other_flop_2(mac_units_4_io_other_flop_2),
    .io_other_flop_3(mac_units_4_io_other_flop_3),
    .io_other_flop_4(mac_units_4_io_other_flop_4),
    .io_flop(mac_units_4_io_flop),
    .io_coef_subch_drc_th(mac_units_4_io_coef_subch_drc_th),
    .io_coef_subch_drc_offset(mac_units_4_io_coef_subch_drc_offset),
    .io_coef_subch_drc_drcen(mac_units_4_io_coef_subch_drc_drcen),
    .io_coef_mainch_ch0_autoloop(mac_units_4_io_coef_mainch_ch0_autoloop),
    .io_coef_mainch_drc_th(mac_units_4_io_coef_mainch_drc_th),
    .io_coef_mainch_drc_offset(mac_units_4_io_coef_mainch_drc_offset),
    .io_coef_mainch_drc_drcen(mac_units_4_io_coef_mainch_drc_drcen)
  );
  CorUnit cor_unit ( // @[dsptop.scala 89:27]
    .clock(cor_unit_clock),
    .reset(cor_unit_reset),
    .io_uopin_ready(cor_unit_io_uopin_ready),
    .io_uopin_valid(cor_unit_io_uopin_valid),
    .io_uopin_bits_cortype(cor_unit_io_uopin_bits_cortype),
    .io_uopin_bits_srcreq_0_valid(cor_unit_io_uopin_bits_srcreq_0_valid),
    .io_uopin_bits_srcreq_0_idx(cor_unit_io_uopin_bits_srcreq_0_idx),
    .io_uopin_bits_srcreq_0_busy(cor_unit_io_uopin_bits_srcreq_0_busy),
    .io_uopin_bits_srcreq_0_wkupidx_0(cor_unit_io_uopin_bits_srcreq_0_wkupidx_0),
    .io_uopin_bits_srcreq_0_wkupidx_1(cor_unit_io_uopin_bits_srcreq_0_wkupidx_1),
    .io_uopin_bits_srcreq_0_wkupidx_2(cor_unit_io_uopin_bits_srcreq_0_wkupidx_2),
    .io_uopin_bits_srcreq_0_wkupidx_3(cor_unit_io_uopin_bits_srcreq_0_wkupidx_3),
    .io_uopin_bits_srcreq_0_wkupidx_4(cor_unit_io_uopin_bits_srcreq_0_wkupidx_4),
    .io_uopin_bits_srcreq_0_wkupidx_5(cor_unit_io_uopin_bits_srcreq_0_wkupidx_5),
    .io_uopin_bits_srcreq_1_valid(cor_unit_io_uopin_bits_srcreq_1_valid),
    .io_uopin_bits_srcreq_1_idx(cor_unit_io_uopin_bits_srcreq_1_idx),
    .io_uopin_bits_srcreq_1_busy(cor_unit_io_uopin_bits_srcreq_1_busy),
    .io_uopin_bits_srcreq_1_wkupidx_0(cor_unit_io_uopin_bits_srcreq_1_wkupidx_0),
    .io_uopin_bits_srcreq_1_wkupidx_1(cor_unit_io_uopin_bits_srcreq_1_wkupidx_1),
    .io_uopin_bits_srcreq_1_wkupidx_2(cor_unit_io_uopin_bits_srcreq_1_wkupidx_2),
    .io_uopin_bits_srcreq_1_wkupidx_3(cor_unit_io_uopin_bits_srcreq_1_wkupidx_3),
    .io_uopin_bits_srcreq_1_wkupidx_4(cor_unit_io_uopin_bits_srcreq_1_wkupidx_4),
    .io_uopin_bits_srcreq_1_wkupidx_5(cor_unit_io_uopin_bits_srcreq_1_wkupidx_5),
    .io_uopin_bits_wbvld(cor_unit_io_uopin_bits_wbvld),
    .io_uopin_bits_wbreq(cor_unit_io_uopin_bits_wbreq),
    .io_uopin_bits_waridx_0(cor_unit_io_uopin_bits_waridx_0),
    .io_uopin_bits_waridx_1(cor_unit_io_uopin_bits_waridx_1),
    .io_uopin_bits_waridx_2(cor_unit_io_uopin_bits_waridx_2),
    .io_uopin_bits_waridx_3(cor_unit_io_uopin_bits_waridx_3),
    .io_uopin_bits_waridx_4(cor_unit_io_uopin_bits_waridx_4),
    .io_uopin_bits_wawidx_0(cor_unit_io_uopin_bits_wawidx_0),
    .io_uopin_bits_wawidx_1(cor_unit_io_uopin_bits_wawidx_1),
    .io_uopin_bits_wawidx_2(cor_unit_io_uopin_bits_wawidx_2),
    .io_uopin_bits_wawidx_3(cor_unit_io_uopin_bits_wawidx_3),
    .io_uopin_bits_wawidx_4(cor_unit_io_uopin_bits_wawidx_4),
    .io_rfreq_0_req_idx(cor_unit_io_rfreq_0_req_idx),
    .io_rfreq_0_resp(cor_unit_io_rfreq_0_resp),
    .io_rfreq_1_req_idx(cor_unit_io_rfreq_1_req_idx),
    .io_rfreq_1_resp(cor_unit_io_rfreq_1_resp),
    .io_wbreq_wdata2(cor_unit_io_wbreq_wdata2),
    .io_wbreq_vld(cor_unit_io_wbreq_vld),
    .io_wbreq_gregidx(cor_unit_io_wbreq_gregidx),
    .io_empty(cor_unit_io_empty),
    .io_fwd_wkup_valid(cor_unit_io_fwd_wkup_valid),
    .io_fwd_wkup_bits(cor_unit_io_fwd_wkup_bits),
    .io_raw_wkup_0_valid(cor_unit_io_raw_wkup_0_valid),
    .io_raw_wkup_0_bits(cor_unit_io_raw_wkup_0_bits),
    .io_raw_wkup_1_valid(cor_unit_io_raw_wkup_1_valid),
    .io_raw_wkup_1_bits(cor_unit_io_raw_wkup_1_bits),
    .io_raw_wkup_2_valid(cor_unit_io_raw_wkup_2_valid),
    .io_raw_wkup_2_bits(cor_unit_io_raw_wkup_2_bits),
    .io_raw_wkup_3_valid(cor_unit_io_raw_wkup_3_valid),
    .io_raw_wkup_3_bits(cor_unit_io_raw_wkup_3_bits),
    .io_raw_wkup_4_valid(cor_unit_io_raw_wkup_4_valid),
    .io_raw_wkup_4_bits(cor_unit_io_raw_wkup_4_bits),
    .io_raw_wkup_5_valid(cor_unit_io_raw_wkup_5_valid),
    .io_raw_wkup_5_bits(cor_unit_io_raw_wkup_5_bits),
    .io_wbcheck_valid(cor_unit_io_wbcheck_valid),
    .io_wbcheck_bits(cor_unit_io_wbcheck_bits),
    .io_r_check_0_valid(cor_unit_io_r_check_0_valid),
    .io_r_check_0_bits(cor_unit_io_r_check_0_bits),
    .io_r_check_1_valid(cor_unit_io_r_check_1_valid),
    .io_r_check_1_bits(cor_unit_io_r_check_1_bits),
    .io_other_flop_0(cor_unit_io_other_flop_0),
    .io_other_flop_1(cor_unit_io_other_flop_1),
    .io_other_flop_2(cor_unit_io_other_flop_2),
    .io_other_flop_3(cor_unit_io_other_flop_3),
    .io_other_flop_4(cor_unit_io_other_flop_4),
    .io_flop(cor_unit_io_flop)
  );
  assign io_din_ready = decode_unit_io_din_ready; // @[dsptop.scala 163:16]
  assign io_dout_valid = decode_unit_io_dout_valid; // @[dsptop.scala 167:17]
  assign io_dout_bits_0 = decode_unit_io_dout_bits_0; // @[dsptop.scala 166:16]
  assign io_dout_bits_1 = decode_unit_io_dout_bits_1; // @[dsptop.scala 166:16]
  assign decode_unit_clock = clock;
  assign decode_unit_reset = reset;
  assign decode_unit_io_din_valid = io_din_valid; // @[dsptop.scala 161:28]
  assign decode_unit_io_din_bits_0 = io_din_bits_0; // @[dsptop.scala 162:27]
  assign decode_unit_io_din_bits_1 = io_din_bits_1; // @[dsptop.scala 162:27]
  assign decode_unit_io_dout_ready = io_dout_ready; // @[dsptop.scala 165:29]
  assign decode_unit_io_macuio_0_ready = mac_units_0_io_uopin_ready; // @[dsptop.scala 171:27]
  assign decode_unit_io_macuio_1_ready = mac_units_1_io_uopin_ready; // @[dsptop.scala 171:27]
  assign decode_unit_io_macuio_2_ready = mac_units_2_io_uopin_ready; // @[dsptop.scala 171:27]
  assign decode_unit_io_macuio_3_ready = mac_units_3_io_uopin_ready; // @[dsptop.scala 171:27]
  assign decode_unit_io_macuio_4_ready = mac_units_4_io_uopin_ready; // @[dsptop.scala 171:27]
  assign decode_unit_io_wd_check_0_valid = mac_units_0_io_wbcheck_valid; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_0_bits = mac_units_0_io_wbcheck_bits; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_1_valid = mac_units_1_io_wbcheck_valid; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_1_bits = mac_units_1_io_wbcheck_bits; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_2_valid = mac_units_2_io_wbcheck_valid; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_2_bits = mac_units_2_io_wbcheck_bits; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_3_valid = mac_units_3_io_wbcheck_valid; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_3_bits = mac_units_3_io_wbcheck_bits; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_4_valid = mac_units_4_io_wbcheck_valid; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_4_bits = mac_units_4_io_wbcheck_bits; // @[dsptop.scala 172:32]
  assign decode_unit_io_wd_check_5_valid = cor_unit_io_wbcheck_valid; // @[dsptop.scala 181:37]
  assign decode_unit_io_wd_check_5_bits = cor_unit_io_wbcheck_bits; // @[dsptop.scala 181:37]
  assign decode_unit_io_mac_r_check_0_0_valid = mac_units_0_io_r_check_0_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_0_bits = mac_units_0_io_r_check_0_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_1_valid = mac_units_0_io_r_check_1_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_1_bits = mac_units_0_io_r_check_1_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_2_valid = mac_units_0_io_r_check_2_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_2_bits = mac_units_0_io_r_check_2_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_3_valid = mac_units_0_io_r_check_3_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_3_bits = mac_units_0_io_r_check_3_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_4_valid = mac_units_0_io_r_check_4_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_4_bits = mac_units_0_io_r_check_4_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_5_valid = mac_units_0_io_r_check_5_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_0_5_bits = mac_units_0_io_r_check_5_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_0_valid = mac_units_1_io_r_check_0_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_0_bits = mac_units_1_io_r_check_0_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_1_valid = mac_units_1_io_r_check_1_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_1_bits = mac_units_1_io_r_check_1_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_2_valid = mac_units_1_io_r_check_2_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_2_bits = mac_units_1_io_r_check_2_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_3_valid = mac_units_1_io_r_check_3_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_3_bits = mac_units_1_io_r_check_3_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_4_valid = mac_units_1_io_r_check_4_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_4_bits = mac_units_1_io_r_check_4_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_5_valid = mac_units_1_io_r_check_5_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_1_5_bits = mac_units_1_io_r_check_5_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_0_valid = mac_units_2_io_r_check_0_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_0_bits = mac_units_2_io_r_check_0_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_1_valid = mac_units_2_io_r_check_1_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_1_bits = mac_units_2_io_r_check_1_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_2_valid = mac_units_2_io_r_check_2_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_2_bits = mac_units_2_io_r_check_2_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_3_valid = mac_units_2_io_r_check_3_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_3_bits = mac_units_2_io_r_check_3_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_4_valid = mac_units_2_io_r_check_4_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_4_bits = mac_units_2_io_r_check_4_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_5_valid = mac_units_2_io_r_check_5_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_2_5_bits = mac_units_2_io_r_check_5_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_0_valid = mac_units_3_io_r_check_0_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_0_bits = mac_units_3_io_r_check_0_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_1_valid = mac_units_3_io_r_check_1_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_1_bits = mac_units_3_io_r_check_1_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_2_valid = mac_units_3_io_r_check_2_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_2_bits = mac_units_3_io_r_check_2_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_3_valid = mac_units_3_io_r_check_3_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_3_bits = mac_units_3_io_r_check_3_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_4_valid = mac_units_3_io_r_check_4_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_4_bits = mac_units_3_io_r_check_4_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_5_valid = mac_units_3_io_r_check_5_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_3_5_bits = mac_units_3_io_r_check_5_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_0_valid = mac_units_4_io_r_check_0_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_0_bits = mac_units_4_io_r_check_0_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_1_valid = mac_units_4_io_r_check_1_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_1_bits = mac_units_4_io_r_check_1_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_2_valid = mac_units_4_io_r_check_2_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_2_bits = mac_units_4_io_r_check_2_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_3_valid = mac_units_4_io_r_check_3_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_3_bits = mac_units_4_io_r_check_3_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_4_valid = mac_units_4_io_r_check_4_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_4_bits = mac_units_4_io_r_check_4_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_5_valid = mac_units_4_io_r_check_5_valid; // @[dsptop.scala 173:35]
  assign decode_unit_io_mac_r_check_4_5_bits = mac_units_4_io_r_check_5_bits; // @[dsptop.scala 173:35]
  assign decode_unit_io_cor_r_check_0_valid = cor_unit_io_r_check_0_valid; // @[dsptop.scala 182:30]
  assign decode_unit_io_cor_r_check_0_bits = cor_unit_io_r_check_0_bits; // @[dsptop.scala 182:30]
  assign decode_unit_io_cor_r_check_1_valid = cor_unit_io_r_check_1_valid; // @[dsptop.scala 182:30]
  assign decode_unit_io_cor_r_check_1_bits = cor_unit_io_r_check_1_bits; // @[dsptop.scala 182:30]
  assign decode_unit_io_exuempty_0 = mac_units_0_io_empty; // @[dsptop.scala 174:32]
  assign decode_unit_io_exuempty_1 = mac_units_1_io_empty; // @[dsptop.scala 174:32]
  assign decode_unit_io_exuempty_2 = mac_units_2_io_empty; // @[dsptop.scala 174:32]
  assign decode_unit_io_exuempty_3 = mac_units_3_io_empty; // @[dsptop.scala 174:32]
  assign decode_unit_io_exuempty_4 = mac_units_4_io_empty; // @[dsptop.scala 174:32]
  assign decode_unit_io_exuempty_5 = cor_unit_io_empty; // @[dsptop.scala 183:37]
  assign decode_unit_io_coruio_ready = cor_unit_io_uopin_ready; // @[dsptop.scala 180:21]
  assign decode_unit_io_readrf_0 = reg_file_io_dec_rd_0; // @[dsptop.scala 177:25]
  assign decode_unit_io_readrf_1 = reg_file_io_dec_rd_1; // @[dsptop.scala 177:25]
  assign decode_unit_io_coef_in_mainch_ch0_inputsel = io_coefin_regmap_mainch_ch1_din_sel; // @[dsptop.scala 90:25 dsptop.scala 111:28]
  assign decode_unit_io_coef_in_mainch_ch1_inputsel = io_coefin_regmap_mainch_ch2_din_sel; // @[dsptop.scala 90:25 dsptop.scala 129:28]
  assign reg_file_clock = clock;
  assign reg_file_reset = reset;
  assign reg_file_io_exe_rd_0_req_isgroup = mac_units_0_io_rfreq_0_req_isgroup; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_0_req_iscoef = mac_units_0_io_rfreq_0_req_iscoef; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_0_req_idx = mac_units_0_io_rfreq_0_req_idx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_0_req_gidx = mac_units_0_io_rfreq_0_req_gidx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_1_req_isgroup = mac_units_0_io_rfreq_1_req_isgroup; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_1_req_iscoef = mac_units_0_io_rfreq_1_req_iscoef; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_1_req_idx = mac_units_0_io_rfreq_1_req_idx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_1_req_gidx = mac_units_0_io_rfreq_1_req_gidx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_1_req_sel = mac_units_0_io_rfreq_1_req_sel; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_2_req_isgroup = mac_units_1_io_rfreq_0_req_isgroup; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_2_req_iscoef = mac_units_1_io_rfreq_0_req_iscoef; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_2_req_idx = mac_units_1_io_rfreq_0_req_idx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_2_req_gidx = mac_units_1_io_rfreq_0_req_gidx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_3_req_isgroup = mac_units_1_io_rfreq_1_req_isgroup; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_3_req_iscoef = mac_units_1_io_rfreq_1_req_iscoef; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_3_req_idx = mac_units_1_io_rfreq_1_req_idx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_3_req_gidx = mac_units_1_io_rfreq_1_req_gidx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_3_req_sel = mac_units_1_io_rfreq_1_req_sel; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_4_req_isgroup = mac_units_2_io_rfreq_0_req_isgroup; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_4_req_iscoef = mac_units_2_io_rfreq_0_req_iscoef; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_4_req_idx = mac_units_2_io_rfreq_0_req_idx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_4_req_gidx = mac_units_2_io_rfreq_0_req_gidx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_5_req_isgroup = mac_units_2_io_rfreq_1_req_isgroup; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_5_req_iscoef = mac_units_2_io_rfreq_1_req_iscoef; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_5_req_idx = mac_units_2_io_rfreq_1_req_idx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_5_req_gidx = mac_units_2_io_rfreq_1_req_gidx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_5_req_sel = mac_units_2_io_rfreq_1_req_sel; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_6_req_isgroup = mac_units_3_io_rfreq_0_req_isgroup; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_6_req_iscoef = mac_units_3_io_rfreq_0_req_iscoef; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_6_req_idx = mac_units_3_io_rfreq_0_req_idx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_6_req_gidx = mac_units_3_io_rfreq_0_req_gidx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_7_req_isgroup = mac_units_3_io_rfreq_1_req_isgroup; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_7_req_iscoef = mac_units_3_io_rfreq_1_req_iscoef; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_7_req_idx = mac_units_3_io_rfreq_1_req_idx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_7_req_gidx = mac_units_3_io_rfreq_1_req_gidx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_7_req_sel = mac_units_3_io_rfreq_1_req_sel; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_8_req_isgroup = mac_units_4_io_rfreq_0_req_isgroup; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_8_req_iscoef = mac_units_4_io_rfreq_0_req_iscoef; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_8_req_idx = mac_units_4_io_rfreq_0_req_idx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_8_req_gidx = mac_units_4_io_rfreq_0_req_gidx; // @[dsptop.scala 192:31]
  assign reg_file_io_exe_rd_9_req_isgroup = mac_units_4_io_rfreq_1_req_isgroup; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_9_req_iscoef = mac_units_4_io_rfreq_1_req_iscoef; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_9_req_idx = mac_units_4_io_rfreq_1_req_idx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_9_req_gidx = mac_units_4_io_rfreq_1_req_gidx; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_9_req_sel = mac_units_4_io_rfreq_1_req_sel; // @[dsptop.scala 193:35]
  assign reg_file_io_exe_rd_10_req_idx = cor_unit_io_rfreq_0_req_idx; // @[dsptop.scala 197:36]
  assign reg_file_io_exe_rd_11_req_idx = cor_unit_io_rfreq_1_req_idx; // @[dsptop.scala 198:40]
  assign reg_file_io_exe_wb_0_wdata1 = mac_units_0_io_wbreq_wdata1; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_0_wdata2 = mac_units_0_io_wbreq_wdata2; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_0_vld = mac_units_0_io_wbreq_vld; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_0_gregidx = mac_units_0_io_wbreq_gregidx; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_1_wdata1 = mac_units_1_io_wbreq_wdata1; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_1_wdata2 = mac_units_1_io_wbreq_wdata2; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_1_vld = mac_units_1_io_wbreq_vld; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_1_gregidx = mac_units_1_io_wbreq_gregidx; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_2_wdata1 = mac_units_2_io_wbreq_wdata1; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_2_wdata2 = mac_units_2_io_wbreq_wdata2; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_2_vld = mac_units_2_io_wbreq_vld; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_2_gregidx = mac_units_2_io_wbreq_gregidx; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_3_wdata1 = mac_units_3_io_wbreq_wdata1; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_3_wdata2 = mac_units_3_io_wbreq_wdata2; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_3_vld = mac_units_3_io_wbreq_vld; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_3_gregidx = mac_units_3_io_wbreq_gregidx; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_4_wdata1 = mac_units_4_io_wbreq_wdata1; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_4_wdata2 = mac_units_4_io_wbreq_wdata2; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_4_vld = mac_units_4_io_wbreq_vld; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_4_gregidx = mac_units_4_io_wbreq_gregidx; // @[dsptop.scala 191:27]
  assign reg_file_io_exe_wb_5_wdata2 = cor_unit_io_wbreq_wdata2; // @[dsptop.scala 196:32]
  assign reg_file_io_exe_wb_5_vld = cor_unit_io_wbreq_vld; // @[dsptop.scala 196:32]
  assign reg_file_io_exe_wb_5_gregidx = cor_unit_io_wbreq_gregidx; // @[dsptop.scala 196:32]
  assign reg_file_io_dec_wb_valid = decode_unit_io_writerf_valid; // @[dsptop.scala 178:22]
  assign reg_file_io_dec_wb_bits_0 = decode_unit_io_writerf_bits_0; // @[dsptop.scala 178:22]
  assign reg_file_io_dec_wb_bits_1 = decode_unit_io_writerf_bits_1; // @[dsptop.scala 178:22]
  assign reg_file_io_dec_wb_bits_2 = decode_unit_io_writerf_bits_2; // @[dsptop.scala 178:22]
  assign reg_file_io_dec_wb_bits_3 = decode_unit_io_writerf_bits_3; // @[dsptop.scala 178:22]
  assign reg_file_io_coef_in_subch_ch2mix_0 = {coef_subch_ch2mix_0_hi,coef_subch_ch2mix_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2mix_1 = {coef_subch_ch2mix_1_hi,coef_subch_ch2mix_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2mix_2 = {coef_subch_ch2mix_2_hi,coef_subch_ch2mix_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2bq_0_0 = {coef_subch_ch2bq_0_0_hi,coef_subch_ch2bq_0_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2bq_0_1 = {coef_subch_ch2bq_0_1_hi,coef_subch_ch2bq_0_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2bq_0_2 = {coef_subch_ch2bq_0_2_hi,coef_subch_ch2bq_0_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2bq_0_3 = {coef_subch_ch2bq_0_3_hi,coef_subch_ch2bq_0_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2bq_0_4 = {coef_subch_ch2bq_0_4_hi,coef_subch_ch2bq_0_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch2vol = io_coefin_regmap_subch_vol_coef; // @[dsptop.scala 90:25 dsptop.scala 145:21]
  assign reg_file_io_coef_in_subch_ch2volsel = io_coefin_regmap_subch_vol_sel[0]; // @[dsptop.scala 90:25 dsptop.scala 146:24]
  assign reg_file_io_coef_in_subch_ch3sel = io_coefin_regmap_subch_ch4_input_sel; // @[dsptop.scala 90:25 dsptop.scala 153:21]
  assign reg_file_io_coef_in_subch_ch3mix_0 = {coef_subch_ch3mix_0_hi,coef_subch_ch3mix_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3mix_1 = {coef_subch_ch3mix_1_hi,coef_subch_ch3mix_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_0_0 = {coef_subch_ch3bq_0_0_hi,coef_subch_ch3bq_0_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_0_1 = {coef_subch_ch3bq_0_1_hi,coef_subch_ch3bq_0_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_0_2 = {coef_subch_ch3bq_0_2_hi,coef_subch_ch3bq_0_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_0_3 = {coef_subch_ch3bq_0_3_hi,coef_subch_ch3bq_0_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_0_4 = {coef_subch_ch3bq_0_4_hi,coef_subch_ch3bq_0_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_1_0 = {coef_subch_ch3bq_1_0_hi,coef_subch_ch3bq_1_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_1_1 = {coef_subch_ch3bq_1_1_hi,coef_subch_ch3bq_1_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_1_2 = {coef_subch_ch3bq_1_2_hi,coef_subch_ch3bq_1_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_1_3 = {coef_subch_ch3bq_1_3_hi,coef_subch_ch3bq_1_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3bq_1_4 = {coef_subch_ch3bq_1_4_hi,coef_subch_ch3bq_1_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_ch3vol = io_coefin_regmap_subch_vol_coef; // @[dsptop.scala 90:25 dsptop.scala 151:21]
  assign reg_file_io_coef_in_subch_ch3volsel = io_coefin_regmap_subch_vol_sel[0]; // @[dsptop.scala 90:25 dsptop.scala 152:24]
  assign reg_file_io_coef_in_subch_drc_pow_0 = {coef_subch_drc_pow_0_hi,coef_subch_drc_pow_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_drc_pow_1 = {coef_subch_drc_pow_1_hi,coef_subch_drc_pow_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_drc_smooth_0 = {coef_subch_drc_smooth_0_hi,coef_subch_drc_smooth_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_drc_smooth_1 = {coef_subch_drc_smooth_1_hi,coef_subch_drc_smooth_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_drc_smooth_2 = {coef_subch_drc_smooth_2_hi,coef_subch_drc_smooth_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_drc_smooth_3 = {coef_subch_drc_smooth_3_hi,coef_subch_drc_smooth_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_subch_drc_ratio = {coef_subch_drc_ratio_hi,coef_subch_drc_ratio_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_0_0 = {coef_mainch_ch0_bqcoef_0_0_hi,coef_mainch_ch0_bqcoef_0_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_0_1 = {coef_mainch_ch0_bqcoef_0_1_hi,coef_mainch_ch0_bqcoef_0_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_0_2 = {coef_mainch_ch0_bqcoef_0_2_hi,coef_mainch_ch0_bqcoef_0_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_0_3 = {coef_mainch_ch0_bqcoef_0_3_hi,coef_mainch_ch0_bqcoef_0_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_0_4 = {coef_mainch_ch0_bqcoef_0_4_hi,coef_mainch_ch0_bqcoef_0_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_1_0 = {coef_mainch_ch0_bqcoef_1_0_hi,coef_mainch_ch0_bqcoef_1_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_1_1 = {coef_mainch_ch0_bqcoef_1_1_hi,coef_mainch_ch0_bqcoef_1_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_1_2 = {coef_mainch_ch0_bqcoef_1_2_hi,coef_mainch_ch0_bqcoef_1_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_1_3 = {coef_mainch_ch0_bqcoef_1_3_hi,coef_mainch_ch0_bqcoef_1_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_1_4 = {coef_mainch_ch0_bqcoef_1_4_hi,coef_mainch_ch0_bqcoef_1_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_2_0 = {coef_mainch_ch0_bqcoef_2_0_hi,coef_mainch_ch0_bqcoef_2_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_2_1 = {coef_mainch_ch0_bqcoef_2_1_hi,coef_mainch_ch0_bqcoef_2_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_2_2 = {coef_mainch_ch0_bqcoef_2_2_hi,coef_mainch_ch0_bqcoef_2_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_2_3 = {coef_mainch_ch0_bqcoef_2_3_hi,coef_mainch_ch0_bqcoef_2_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_2_4 = {coef_mainch_ch0_bqcoef_2_4_hi,coef_mainch_ch0_bqcoef_2_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_3_0 = {coef_mainch_ch0_bqcoef_3_0_hi,coef_mainch_ch0_bqcoef_3_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_3_1 = {coef_mainch_ch0_bqcoef_3_1_hi,coef_mainch_ch0_bqcoef_3_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_3_2 = {coef_mainch_ch0_bqcoef_3_2_hi,coef_mainch_ch0_bqcoef_3_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_3_3 = {coef_mainch_ch0_bqcoef_3_3_hi,coef_mainch_ch0_bqcoef_3_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_3_4 = {coef_mainch_ch0_bqcoef_3_4_hi,coef_mainch_ch0_bqcoef_3_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_4_0 = {coef_mainch_ch0_bqcoef_4_0_hi,coef_mainch_ch0_bqcoef_4_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_4_1 = {coef_mainch_ch0_bqcoef_4_1_hi,coef_mainch_ch0_bqcoef_4_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_4_2 = {coef_mainch_ch0_bqcoef_4_2_hi,coef_mainch_ch0_bqcoef_4_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_4_3 = {coef_mainch_ch0_bqcoef_4_3_hi,coef_mainch_ch0_bqcoef_4_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_4_4 = {coef_mainch_ch0_bqcoef_4_4_hi,coef_mainch_ch0_bqcoef_4_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_5_0 = {coef_mainch_ch0_bqcoef_5_0_hi,coef_mainch_ch0_bqcoef_5_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_5_1 = {coef_mainch_ch0_bqcoef_5_1_hi,coef_mainch_ch0_bqcoef_5_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_5_2 = {coef_mainch_ch0_bqcoef_5_2_hi,coef_mainch_ch0_bqcoef_5_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_5_3 = {coef_mainch_ch0_bqcoef_5_3_hi,coef_mainch_ch0_bqcoef_5_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_5_4 = {coef_mainch_ch0_bqcoef_5_4_hi,coef_mainch_ch0_bqcoef_5_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_6_0 = {coef_mainch_ch0_bqcoef_6_0_hi,coef_mainch_ch0_bqcoef_6_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_6_1 = {coef_mainch_ch0_bqcoef_6_1_hi,coef_mainch_ch0_bqcoef_6_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_6_2 = {coef_mainch_ch0_bqcoef_6_2_hi,coef_mainch_ch0_bqcoef_6_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_6_3 = {coef_mainch_ch0_bqcoef_6_3_hi,coef_mainch_ch0_bqcoef_6_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_6_4 = {coef_mainch_ch0_bqcoef_6_4_hi,coef_mainch_ch0_bqcoef_6_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_7_0 = {coef_mainch_ch0_bqcoef_7_0_hi,coef_mainch_ch0_bqcoef_7_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_7_1 = {coef_mainch_ch0_bqcoef_7_1_hi,coef_mainch_ch0_bqcoef_7_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_7_2 = {coef_mainch_ch0_bqcoef_7_2_hi,coef_mainch_ch0_bqcoef_7_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_7_3 = {coef_mainch_ch0_bqcoef_7_3_hi,coef_mainch_ch0_bqcoef_7_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_7_4 = {coef_mainch_ch0_bqcoef_7_4_hi,coef_mainch_ch0_bqcoef_7_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_8_0 = {coef_mainch_ch0_bqcoef_8_0_hi,coef_mainch_ch0_bqcoef_8_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_8_1 = {coef_mainch_ch0_bqcoef_8_1_hi,coef_mainch_ch0_bqcoef_8_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_8_2 = {coef_mainch_ch0_bqcoef_8_2_hi,coef_mainch_ch0_bqcoef_8_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_8_3 = {coef_mainch_ch0_bqcoef_8_3_hi,coef_mainch_ch0_bqcoef_8_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_bqcoef_8_4 = {coef_mainch_ch0_bqcoef_8_4_hi,coef_mainch_ch0_bqcoef_8_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_inputmix_0_0 = {coef_mainch_ch0_inputmix_0_0_hi,coef_mainch_ch0_inputmix_0_0_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_inputmix_0_1 = {coef_mainch_ch0_inputmix_0_1_hi,coef_mainch_ch0_inputmix_0_1_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_inputmix_1_0 = {coef_mainch_ch0_inputmix_1_0_hi,coef_mainch_ch0_inputmix_1_0_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_inputmix_1_1 = {coef_mainch_ch0_inputmix_1_1_hi,coef_mainch_ch0_inputmix_1_1_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_vol = io_coefin_regmap_mainch_ch1_vol_coef; // @[dsptop.scala 90:25 dsptop.scala 110:23]
  assign reg_file_io_coef_in_mainch_ch0_outputmix_0 = {coef_mainch_ch0_outputmix_0_hi,coef_mainch_ch0_outputmix_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_outputmix_1 = {coef_mainch_ch0_outputmix_1_hi,coef_mainch_ch0_outputmix_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_outputmix_2 = {coef_mainch_ch0_outputmix_2_hi,coef_mainch_ch0_outputmix_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch0_prescale = io_coefin_regmap_mainch_pre_scale; // @[dsptop.scala 90:25 dsptop.scala 112:28]
  assign reg_file_io_coef_in_mainch_ch0_postscale = {coef_mainch_ch0_postscale_hi,coef_mainch_ch0_postscale_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_0_0 = {coef_mainch_ch1_bqcoef_0_0_hi,coef_mainch_ch1_bqcoef_0_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_0_1 = {coef_mainch_ch1_bqcoef_0_1_hi,coef_mainch_ch1_bqcoef_0_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_0_2 = {coef_mainch_ch1_bqcoef_0_2_hi,coef_mainch_ch1_bqcoef_0_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_0_3 = {coef_mainch_ch1_bqcoef_0_3_hi,coef_mainch_ch1_bqcoef_0_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_0_4 = {coef_mainch_ch1_bqcoef_0_4_hi,coef_mainch_ch1_bqcoef_0_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_1_0 = {coef_mainch_ch1_bqcoef_1_0_hi,coef_mainch_ch1_bqcoef_1_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_1_1 = {coef_mainch_ch1_bqcoef_1_1_hi,coef_mainch_ch1_bqcoef_1_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_1_2 = {coef_mainch_ch1_bqcoef_1_2_hi,coef_mainch_ch1_bqcoef_1_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_1_3 = {coef_mainch_ch1_bqcoef_1_3_hi,coef_mainch_ch1_bqcoef_1_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_1_4 = {coef_mainch_ch1_bqcoef_1_4_hi,coef_mainch_ch1_bqcoef_1_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_2_0 = {coef_mainch_ch1_bqcoef_2_0_hi,coef_mainch_ch1_bqcoef_2_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_2_1 = {coef_mainch_ch1_bqcoef_2_1_hi,coef_mainch_ch1_bqcoef_2_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_2_2 = {coef_mainch_ch1_bqcoef_2_2_hi,coef_mainch_ch1_bqcoef_2_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_2_3 = {coef_mainch_ch1_bqcoef_2_3_hi,coef_mainch_ch1_bqcoef_2_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_2_4 = {coef_mainch_ch1_bqcoef_2_4_hi,coef_mainch_ch1_bqcoef_2_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_3_0 = {coef_mainch_ch1_bqcoef_3_0_hi,coef_mainch_ch1_bqcoef_3_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_3_1 = {coef_mainch_ch1_bqcoef_3_1_hi,coef_mainch_ch1_bqcoef_3_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_3_2 = {coef_mainch_ch1_bqcoef_3_2_hi,coef_mainch_ch1_bqcoef_3_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_3_3 = {coef_mainch_ch1_bqcoef_3_3_hi,coef_mainch_ch1_bqcoef_3_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_3_4 = {coef_mainch_ch1_bqcoef_3_4_hi,coef_mainch_ch1_bqcoef_3_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_4_0 = {coef_mainch_ch1_bqcoef_4_0_hi,coef_mainch_ch1_bqcoef_4_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_4_1 = {coef_mainch_ch1_bqcoef_4_1_hi,coef_mainch_ch1_bqcoef_4_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_4_2 = {coef_mainch_ch1_bqcoef_4_2_hi,coef_mainch_ch1_bqcoef_4_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_4_3 = {coef_mainch_ch1_bqcoef_4_3_hi,coef_mainch_ch1_bqcoef_4_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_4_4 = {coef_mainch_ch1_bqcoef_4_4_hi,coef_mainch_ch1_bqcoef_4_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_5_0 = {coef_mainch_ch1_bqcoef_5_0_hi,coef_mainch_ch1_bqcoef_5_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_5_1 = {coef_mainch_ch1_bqcoef_5_1_hi,coef_mainch_ch1_bqcoef_5_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_5_2 = {coef_mainch_ch1_bqcoef_5_2_hi,coef_mainch_ch1_bqcoef_5_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_5_3 = {coef_mainch_ch1_bqcoef_5_3_hi,coef_mainch_ch1_bqcoef_5_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_5_4 = {coef_mainch_ch1_bqcoef_5_4_hi,coef_mainch_ch1_bqcoef_5_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_6_0 = {coef_mainch_ch1_bqcoef_6_0_hi,coef_mainch_ch1_bqcoef_6_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_6_1 = {coef_mainch_ch1_bqcoef_6_1_hi,coef_mainch_ch1_bqcoef_6_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_6_2 = {coef_mainch_ch1_bqcoef_6_2_hi,coef_mainch_ch1_bqcoef_6_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_6_3 = {coef_mainch_ch1_bqcoef_6_3_hi,coef_mainch_ch1_bqcoef_6_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_6_4 = {coef_mainch_ch1_bqcoef_6_4_hi,coef_mainch_ch1_bqcoef_6_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_7_0 = {coef_mainch_ch1_bqcoef_7_0_hi,coef_mainch_ch1_bqcoef_7_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_7_1 = {coef_mainch_ch1_bqcoef_7_1_hi,coef_mainch_ch1_bqcoef_7_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_7_2 = {coef_mainch_ch1_bqcoef_7_2_hi,coef_mainch_ch1_bqcoef_7_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_7_3 = {coef_mainch_ch1_bqcoef_7_3_hi,coef_mainch_ch1_bqcoef_7_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_7_4 = {coef_mainch_ch1_bqcoef_7_4_hi,coef_mainch_ch1_bqcoef_7_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_8_0 = {coef_mainch_ch1_bqcoef_8_0_hi,coef_mainch_ch1_bqcoef_8_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_8_1 = {coef_mainch_ch1_bqcoef_8_1_hi,coef_mainch_ch1_bqcoef_8_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_8_2 = {coef_mainch_ch1_bqcoef_8_2_hi,coef_mainch_ch1_bqcoef_8_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_8_3 = {coef_mainch_ch1_bqcoef_8_3_hi,coef_mainch_ch1_bqcoef_8_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_bqcoef_8_4 = {coef_mainch_ch1_bqcoef_8_4_hi,coef_mainch_ch1_bqcoef_8_4_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_inputmix_0_0 = {coef_mainch_ch1_inputmix_0_0_hi,coef_mainch_ch1_inputmix_0_0_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_inputmix_0_1 = {coef_mainch_ch1_inputmix_0_1_hi,coef_mainch_ch1_inputmix_0_1_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_inputmix_1_0 = {coef_mainch_ch1_inputmix_1_0_hi,coef_mainch_ch1_inputmix_1_0_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_inputmix_1_1 = {coef_mainch_ch1_inputmix_1_1_hi,coef_mainch_ch1_inputmix_1_1_lo}
    ; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_vol = io_coefin_regmap_mainch_ch2_vol_coef; // @[dsptop.scala 90:25 dsptop.scala 128:23]
  assign reg_file_io_coef_in_mainch_ch1_outputmix_0 = {coef_mainch_ch1_outputmix_0_hi,coef_mainch_ch1_outputmix_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_outputmix_1 = {coef_mainch_ch1_outputmix_1_hi,coef_mainch_ch1_outputmix_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_ch1_outputmix_2 = {coef_mainch_ch1_outputmix_2_hi,coef_mainch_ch1_outputmix_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_pow_0 = {coef_mainch_drc_pow_0_hi,coef_mainch_drc_pow_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_pow_1 = {coef_mainch_drc_pow_1_hi,coef_mainch_drc_pow_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_smooth_0 = {coef_mainch_drc_smooth_0_hi,coef_mainch_drc_smooth_0_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_smooth_1 = {coef_mainch_drc_smooth_1_hi,coef_mainch_drc_smooth_1_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_smooth_2 = {coef_mainch_drc_smooth_2_hi,coef_mainch_drc_smooth_2_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_smooth_3 = {coef_mainch_drc_smooth_3_hi,coef_mainch_drc_smooth_3_lo}; // @[Cat.scala 30:58]
  assign reg_file_io_coef_in_mainch_drc_ratio = {coef_mainch_drc_ratio_hi,coef_mainch_drc_ratio_lo}; // @[Cat.scala 30:58]
  assign mac_units_0_clock = clock;
  assign mac_units_0_reset = reset;
  assign mac_units_0_io_uopin_valid = decode_unit_io_macuio_0_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_vlen = decode_unit_io_macuio_0_bits_vlen; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_select = decode_unit_io_macuio_0_bits_select; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_drc = decode_unit_io_macuio_0_bits_drc; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_pow = decode_unit_io_macuio_0_bits_pow; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_loop = decode_unit_io_macuio_0_bits_loop; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_drcgain = decode_unit_io_macuio_0_bits_drcgain; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_drcnum = decode_unit_io_macuio_0_bits_drcnum; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_valid = decode_unit_io_macuio_0_bits_srcreq_0_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_isgroup = decode_unit_io_macuio_0_bits_srcreq_0_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_iscoef = decode_unit_io_macuio_0_bits_srcreq_0_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_idx = decode_unit_io_macuio_0_bits_srcreq_0_idx; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_busy = decode_unit_io_macuio_0_bits_srcreq_0_busy; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_wkupidx_0 = decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_wkupidx_1 = decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_wkupidx_2 = decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_wkupidx_3 = decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_wkupidx_4 = decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_0_wkupidx_5 = decode_unit_io_macuio_0_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_valid = decode_unit_io_macuio_0_bits_srcreq_1_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_isgroup = decode_unit_io_macuio_0_bits_srcreq_1_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_iscoef = decode_unit_io_macuio_0_bits_srcreq_1_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_idx = decode_unit_io_macuio_0_bits_srcreq_1_idx; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_busy = decode_unit_io_macuio_0_bits_srcreq_1_busy; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_wkupidx_0 = decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_wkupidx_1 = decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_wkupidx_2 = decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_wkupidx_3 = decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_wkupidx_4 = decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_1_wkupidx_5 = decode_unit_io_macuio_0_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_valid = decode_unit_io_macuio_0_bits_srcreq_2_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_isgroup = decode_unit_io_macuio_0_bits_srcreq_2_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_iscoef = decode_unit_io_macuio_0_bits_srcreq_2_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_idx = decode_unit_io_macuio_0_bits_srcreq_2_idx; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_busy = decode_unit_io_macuio_0_bits_srcreq_2_busy; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_wkupidx_0 = decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_wkupidx_1 = decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_wkupidx_2 = decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_wkupidx_3 = decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_wkupidx_4 = decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_2_wkupidx_5 = decode_unit_io_macuio_0_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_valid = decode_unit_io_macuio_0_bits_srcreq_3_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_isgroup = decode_unit_io_macuio_0_bits_srcreq_3_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_iscoef = decode_unit_io_macuio_0_bits_srcreq_3_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_idx = decode_unit_io_macuio_0_bits_srcreq_3_idx; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_busy = decode_unit_io_macuio_0_bits_srcreq_3_busy; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_wkupidx_0 = decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_wkupidx_1 = decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_wkupidx_2 = decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_wkupidx_3 = decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_wkupidx_4 = decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_3_wkupidx_5 = decode_unit_io_macuio_0_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_valid = decode_unit_io_macuio_0_bits_srcreq_4_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_isgroup = decode_unit_io_macuio_0_bits_srcreq_4_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_iscoef = decode_unit_io_macuio_0_bits_srcreq_4_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_idx = decode_unit_io_macuio_0_bits_srcreq_4_idx; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_busy = decode_unit_io_macuio_0_bits_srcreq_4_busy; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_wkupidx_0 = decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_wkupidx_1 = decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_wkupidx_2 = decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_wkupidx_3 = decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_wkupidx_4 = decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_4_wkupidx_5 = decode_unit_io_macuio_0_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_valid = decode_unit_io_macuio_0_bits_srcreq_5_valid; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_isgroup = decode_unit_io_macuio_0_bits_srcreq_5_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_iscoef = decode_unit_io_macuio_0_bits_srcreq_5_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_idx = decode_unit_io_macuio_0_bits_srcreq_5_idx; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_busy = decode_unit_io_macuio_0_bits_srcreq_5_busy; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_wkupidx_0 = decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_wkupidx_1 = decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_wkupidx_2 = decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_wkupidx_3 = decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_wkupidx_4 = decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_srcreq_5_wkupidx_5 = decode_unit_io_macuio_0_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wbvld = decode_unit_io_macuio_0_bits_wbvld; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wbreq = decode_unit_io_macuio_0_bits_wbreq; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_waridx_0 = decode_unit_io_macuio_0_bits_waridx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_waridx_1 = decode_unit_io_macuio_0_bits_waridx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_waridx_2 = decode_unit_io_macuio_0_bits_waridx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_waridx_3 = decode_unit_io_macuio_0_bits_waridx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_waridx_4 = decode_unit_io_macuio_0_bits_waridx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wawidx_0 = decode_unit_io_macuio_0_bits_wawidx_0; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wawidx_1 = decode_unit_io_macuio_0_bits_wawidx_1; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wawidx_2 = decode_unit_io_macuio_0_bits_wawidx_2; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wawidx_3 = decode_unit_io_macuio_0_bits_wawidx_3; // @[dsptop.scala 171:27]
  assign mac_units_0_io_uopin_bits_wawidx_4 = decode_unit_io_macuio_0_bits_wawidx_4; // @[dsptop.scala 171:27]
  assign mac_units_0_io_rfreq_0_resp = reg_file_io_exe_rd_0_resp; // @[dsptop.scala 192:31]
  assign mac_units_0_io_rfreq_1_resp = reg_file_io_exe_rd_1_resp; // @[dsptop.scala 193:35]
  assign mac_units_0_io_raw_wkup_0_valid = mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_0_bits = mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_1_valid = mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_1_bits = mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_2_valid = mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_2_bits = mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_3_valid = mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_3_bits = mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_4_valid = mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_4_bits = mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_0_io_raw_wkup_5_valid = cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_0_io_raw_wkup_5_bits = cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_0_io_other_flop_0 = mac_units_1_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_0_io_other_flop_1 = mac_units_2_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_0_io_other_flop_2 = mac_units_3_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_0_io_other_flop_3 = mac_units_4_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_0_io_other_flop_4 = cor_unit_io_flop; // @[dsptop.scala 205:25 dsptop.scala 216:22]
  assign mac_units_0_io_coef_subch_drc_th = io_coefin_regmap_subch_drc2_coef[95:64]; // @[dsptop.scala 105:56]
  assign mac_units_0_io_coef_subch_drc_offset = {coef_subch_drc_offset_hi,coef_subch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_0_io_coef_subch_drc_drcen = io_coefin_regmap_subch_drc2_en; // @[dsptop.scala 90:25 dsptop.scala 102:24]
  assign mac_units_0_io_coef_mainch_ch0_autoloop = io_coefin_regmap_mainch_alp_en; // @[dsptop.scala 90:25 dsptop.scala 109:28]
  assign mac_units_0_io_coef_mainch_drc_th = io_coefin_regmap_mainch_drc1_coef[95:64]; // @[dsptop.scala 98:58]
  assign mac_units_0_io_coef_mainch_drc_offset = {coef_mainch_drc_offset_hi,coef_mainch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_0_io_coef_mainch_drc_drcen = io_coefin_regmap_mainch_drc1_en; // @[dsptop.scala 90:25 dsptop.scala 95:25]
  assign mac_units_1_clock = clock;
  assign mac_units_1_reset = reset;
  assign mac_units_1_io_uopin_valid = decode_unit_io_macuio_1_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_vlen = decode_unit_io_macuio_1_bits_vlen; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_select = decode_unit_io_macuio_1_bits_select; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_drc = decode_unit_io_macuio_1_bits_drc; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_pow = decode_unit_io_macuio_1_bits_pow; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_loop = decode_unit_io_macuio_1_bits_loop; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_drcgain = decode_unit_io_macuio_1_bits_drcgain; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_drcnum = decode_unit_io_macuio_1_bits_drcnum; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_valid = decode_unit_io_macuio_1_bits_srcreq_0_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_isgroup = decode_unit_io_macuio_1_bits_srcreq_0_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_iscoef = decode_unit_io_macuio_1_bits_srcreq_0_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_idx = decode_unit_io_macuio_1_bits_srcreq_0_idx; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_busy = decode_unit_io_macuio_1_bits_srcreq_0_busy; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_wkupidx_0 = decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_wkupidx_1 = decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_wkupidx_2 = decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_wkupidx_3 = decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_wkupidx_4 = decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_0_wkupidx_5 = decode_unit_io_macuio_1_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_valid = decode_unit_io_macuio_1_bits_srcreq_1_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_isgroup = decode_unit_io_macuio_1_bits_srcreq_1_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_iscoef = decode_unit_io_macuio_1_bits_srcreq_1_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_idx = decode_unit_io_macuio_1_bits_srcreq_1_idx; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_busy = decode_unit_io_macuio_1_bits_srcreq_1_busy; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_wkupidx_0 = decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_wkupidx_1 = decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_wkupidx_2 = decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_wkupidx_3 = decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_wkupidx_4 = decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_1_wkupidx_5 = decode_unit_io_macuio_1_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_valid = decode_unit_io_macuio_1_bits_srcreq_2_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_isgroup = decode_unit_io_macuio_1_bits_srcreq_2_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_iscoef = decode_unit_io_macuio_1_bits_srcreq_2_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_idx = decode_unit_io_macuio_1_bits_srcreq_2_idx; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_busy = decode_unit_io_macuio_1_bits_srcreq_2_busy; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_wkupidx_0 = decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_wkupidx_1 = decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_wkupidx_2 = decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_wkupidx_3 = decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_wkupidx_4 = decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_2_wkupidx_5 = decode_unit_io_macuio_1_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_valid = decode_unit_io_macuio_1_bits_srcreq_3_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_isgroup = decode_unit_io_macuio_1_bits_srcreq_3_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_iscoef = decode_unit_io_macuio_1_bits_srcreq_3_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_idx = decode_unit_io_macuio_1_bits_srcreq_3_idx; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_busy = decode_unit_io_macuio_1_bits_srcreq_3_busy; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_wkupidx_0 = decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_wkupidx_1 = decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_wkupidx_2 = decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_wkupidx_3 = decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_wkupidx_4 = decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_3_wkupidx_5 = decode_unit_io_macuio_1_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_valid = decode_unit_io_macuio_1_bits_srcreq_4_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_isgroup = decode_unit_io_macuio_1_bits_srcreq_4_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_iscoef = decode_unit_io_macuio_1_bits_srcreq_4_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_idx = decode_unit_io_macuio_1_bits_srcreq_4_idx; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_busy = decode_unit_io_macuio_1_bits_srcreq_4_busy; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_wkupidx_0 = decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_wkupidx_1 = decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_wkupidx_2 = decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_wkupidx_3 = decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_wkupidx_4 = decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_4_wkupidx_5 = decode_unit_io_macuio_1_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_valid = decode_unit_io_macuio_1_bits_srcreq_5_valid; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_isgroup = decode_unit_io_macuio_1_bits_srcreq_5_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_iscoef = decode_unit_io_macuio_1_bits_srcreq_5_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_idx = decode_unit_io_macuio_1_bits_srcreq_5_idx; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_busy = decode_unit_io_macuio_1_bits_srcreq_5_busy; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_wkupidx_0 = decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_wkupidx_1 = decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_wkupidx_2 = decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_wkupidx_3 = decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_wkupidx_4 = decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_srcreq_5_wkupidx_5 = decode_unit_io_macuio_1_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wbvld = decode_unit_io_macuio_1_bits_wbvld; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wbreq = decode_unit_io_macuio_1_bits_wbreq; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_waridx_0 = decode_unit_io_macuio_1_bits_waridx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_waridx_1 = decode_unit_io_macuio_1_bits_waridx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_waridx_2 = decode_unit_io_macuio_1_bits_waridx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_waridx_3 = decode_unit_io_macuio_1_bits_waridx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_waridx_4 = decode_unit_io_macuio_1_bits_waridx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wawidx_0 = decode_unit_io_macuio_1_bits_wawidx_0; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wawidx_1 = decode_unit_io_macuio_1_bits_wawidx_1; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wawidx_2 = decode_unit_io_macuio_1_bits_wawidx_2; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wawidx_3 = decode_unit_io_macuio_1_bits_wawidx_3; // @[dsptop.scala 171:27]
  assign mac_units_1_io_uopin_bits_wawidx_4 = decode_unit_io_macuio_1_bits_wawidx_4; // @[dsptop.scala 171:27]
  assign mac_units_1_io_rfreq_0_resp = reg_file_io_exe_rd_2_resp; // @[dsptop.scala 192:31]
  assign mac_units_1_io_rfreq_1_resp = reg_file_io_exe_rd_3_resp; // @[dsptop.scala 193:35]
  assign mac_units_1_io_raw_wkup_0_valid = mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_0_bits = mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_1_valid = mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_1_bits = mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_2_valid = mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_2_bits = mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_3_valid = mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_3_bits = mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_4_valid = mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_4_bits = mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_1_io_raw_wkup_5_valid = cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_1_io_raw_wkup_5_bits = cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_1_io_other_flop_0 = mac_units_0_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_1_io_other_flop_1 = mac_units_2_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_1_io_other_flop_2 = mac_units_3_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_1_io_other_flop_3 = mac_units_4_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_1_io_other_flop_4 = cor_unit_io_flop; // @[dsptop.scala 205:25 dsptop.scala 216:22]
  assign mac_units_1_io_coef_subch_drc_th = io_coefin_regmap_subch_drc2_coef[95:64]; // @[dsptop.scala 105:56]
  assign mac_units_1_io_coef_subch_drc_offset = {coef_subch_drc_offset_hi,coef_subch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_1_io_coef_subch_drc_drcen = io_coefin_regmap_subch_drc2_en; // @[dsptop.scala 90:25 dsptop.scala 102:24]
  assign mac_units_1_io_coef_mainch_ch0_autoloop = io_coefin_regmap_mainch_alp_en; // @[dsptop.scala 90:25 dsptop.scala 109:28]
  assign mac_units_1_io_coef_mainch_drc_th = io_coefin_regmap_mainch_drc1_coef[95:64]; // @[dsptop.scala 98:58]
  assign mac_units_1_io_coef_mainch_drc_offset = {coef_mainch_drc_offset_hi,coef_mainch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_1_io_coef_mainch_drc_drcen = io_coefin_regmap_mainch_drc1_en; // @[dsptop.scala 90:25 dsptop.scala 95:25]
  assign mac_units_2_clock = clock;
  assign mac_units_2_reset = reset;
  assign mac_units_2_io_uopin_valid = decode_unit_io_macuio_2_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_vlen = decode_unit_io_macuio_2_bits_vlen; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_select = decode_unit_io_macuio_2_bits_select; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_drc = decode_unit_io_macuio_2_bits_drc; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_pow = decode_unit_io_macuio_2_bits_pow; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_loop = decode_unit_io_macuio_2_bits_loop; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_drcgain = decode_unit_io_macuio_2_bits_drcgain; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_drcnum = decode_unit_io_macuio_2_bits_drcnum; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_valid = decode_unit_io_macuio_2_bits_srcreq_0_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_isgroup = decode_unit_io_macuio_2_bits_srcreq_0_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_iscoef = decode_unit_io_macuio_2_bits_srcreq_0_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_idx = decode_unit_io_macuio_2_bits_srcreq_0_idx; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_busy = decode_unit_io_macuio_2_bits_srcreq_0_busy; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_wkupidx_0 = decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_wkupidx_1 = decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_wkupidx_2 = decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_wkupidx_3 = decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_wkupidx_4 = decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_0_wkupidx_5 = decode_unit_io_macuio_2_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_valid = decode_unit_io_macuio_2_bits_srcreq_1_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_isgroup = decode_unit_io_macuio_2_bits_srcreq_1_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_iscoef = decode_unit_io_macuio_2_bits_srcreq_1_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_idx = decode_unit_io_macuio_2_bits_srcreq_1_idx; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_busy = decode_unit_io_macuio_2_bits_srcreq_1_busy; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_wkupidx_0 = decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_wkupidx_1 = decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_wkupidx_2 = decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_wkupidx_3 = decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_wkupidx_4 = decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_1_wkupidx_5 = decode_unit_io_macuio_2_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_valid = decode_unit_io_macuio_2_bits_srcreq_2_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_isgroup = decode_unit_io_macuio_2_bits_srcreq_2_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_iscoef = decode_unit_io_macuio_2_bits_srcreq_2_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_idx = decode_unit_io_macuio_2_bits_srcreq_2_idx; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_busy = decode_unit_io_macuio_2_bits_srcreq_2_busy; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_wkupidx_0 = decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_wkupidx_1 = decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_wkupidx_2 = decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_wkupidx_3 = decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_wkupidx_4 = decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_2_wkupidx_5 = decode_unit_io_macuio_2_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_valid = decode_unit_io_macuio_2_bits_srcreq_3_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_isgroup = decode_unit_io_macuio_2_bits_srcreq_3_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_iscoef = decode_unit_io_macuio_2_bits_srcreq_3_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_idx = decode_unit_io_macuio_2_bits_srcreq_3_idx; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_busy = decode_unit_io_macuio_2_bits_srcreq_3_busy; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_wkupidx_0 = decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_wkupidx_1 = decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_wkupidx_2 = decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_wkupidx_3 = decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_wkupidx_4 = decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_3_wkupidx_5 = decode_unit_io_macuio_2_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_valid = decode_unit_io_macuio_2_bits_srcreq_4_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_isgroup = decode_unit_io_macuio_2_bits_srcreq_4_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_iscoef = decode_unit_io_macuio_2_bits_srcreq_4_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_idx = decode_unit_io_macuio_2_bits_srcreq_4_idx; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_busy = decode_unit_io_macuio_2_bits_srcreq_4_busy; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_wkupidx_0 = decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_wkupidx_1 = decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_wkupidx_2 = decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_wkupidx_3 = decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_wkupidx_4 = decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_4_wkupidx_5 = decode_unit_io_macuio_2_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_valid = decode_unit_io_macuio_2_bits_srcreq_5_valid; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_isgroup = decode_unit_io_macuio_2_bits_srcreq_5_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_iscoef = decode_unit_io_macuio_2_bits_srcreq_5_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_idx = decode_unit_io_macuio_2_bits_srcreq_5_idx; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_busy = decode_unit_io_macuio_2_bits_srcreq_5_busy; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_wkupidx_0 = decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_wkupidx_1 = decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_wkupidx_2 = decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_wkupidx_3 = decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_wkupidx_4 = decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_srcreq_5_wkupidx_5 = decode_unit_io_macuio_2_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wbvld = decode_unit_io_macuio_2_bits_wbvld; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wbreq = decode_unit_io_macuio_2_bits_wbreq; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_waridx_0 = decode_unit_io_macuio_2_bits_waridx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_waridx_1 = decode_unit_io_macuio_2_bits_waridx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_waridx_2 = decode_unit_io_macuio_2_bits_waridx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_waridx_3 = decode_unit_io_macuio_2_bits_waridx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_waridx_4 = decode_unit_io_macuio_2_bits_waridx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wawidx_0 = decode_unit_io_macuio_2_bits_wawidx_0; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wawidx_1 = decode_unit_io_macuio_2_bits_wawidx_1; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wawidx_2 = decode_unit_io_macuio_2_bits_wawidx_2; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wawidx_3 = decode_unit_io_macuio_2_bits_wawidx_3; // @[dsptop.scala 171:27]
  assign mac_units_2_io_uopin_bits_wawidx_4 = decode_unit_io_macuio_2_bits_wawidx_4; // @[dsptop.scala 171:27]
  assign mac_units_2_io_rfreq_0_resp = reg_file_io_exe_rd_4_resp; // @[dsptop.scala 192:31]
  assign mac_units_2_io_rfreq_1_resp = reg_file_io_exe_rd_5_resp; // @[dsptop.scala 193:35]
  assign mac_units_2_io_raw_wkup_0_valid = mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_0_bits = mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_1_valid = mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_1_bits = mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_2_valid = mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_2_bits = mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_3_valid = mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_3_bits = mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_4_valid = mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_4_bits = mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_2_io_raw_wkup_5_valid = cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_2_io_raw_wkup_5_bits = cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_2_io_other_flop_0 = mac_units_0_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_2_io_other_flop_1 = mac_units_1_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_2_io_other_flop_2 = mac_units_3_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_2_io_other_flop_3 = mac_units_4_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_2_io_other_flop_4 = cor_unit_io_flop; // @[dsptop.scala 205:25 dsptop.scala 216:22]
  assign mac_units_2_io_coef_subch_drc_th = io_coefin_regmap_subch_drc2_coef[95:64]; // @[dsptop.scala 105:56]
  assign mac_units_2_io_coef_subch_drc_offset = {coef_subch_drc_offset_hi,coef_subch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_2_io_coef_subch_drc_drcen = io_coefin_regmap_subch_drc2_en; // @[dsptop.scala 90:25 dsptop.scala 102:24]
  assign mac_units_2_io_coef_mainch_ch0_autoloop = io_coefin_regmap_mainch_alp_en; // @[dsptop.scala 90:25 dsptop.scala 109:28]
  assign mac_units_2_io_coef_mainch_drc_th = io_coefin_regmap_mainch_drc1_coef[95:64]; // @[dsptop.scala 98:58]
  assign mac_units_2_io_coef_mainch_drc_offset = {coef_mainch_drc_offset_hi,coef_mainch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_2_io_coef_mainch_drc_drcen = io_coefin_regmap_mainch_drc1_en; // @[dsptop.scala 90:25 dsptop.scala 95:25]
  assign mac_units_3_clock = clock;
  assign mac_units_3_reset = reset;
  assign mac_units_3_io_uopin_valid = decode_unit_io_macuio_3_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_vlen = decode_unit_io_macuio_3_bits_vlen; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_select = decode_unit_io_macuio_3_bits_select; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_drc = decode_unit_io_macuio_3_bits_drc; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_pow = decode_unit_io_macuio_3_bits_pow; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_loop = decode_unit_io_macuio_3_bits_loop; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_drcgain = decode_unit_io_macuio_3_bits_drcgain; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_drcnum = decode_unit_io_macuio_3_bits_drcnum; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_valid = decode_unit_io_macuio_3_bits_srcreq_0_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_isgroup = decode_unit_io_macuio_3_bits_srcreq_0_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_iscoef = decode_unit_io_macuio_3_bits_srcreq_0_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_idx = decode_unit_io_macuio_3_bits_srcreq_0_idx; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_busy = decode_unit_io_macuio_3_bits_srcreq_0_busy; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_wkupidx_0 = decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_wkupidx_1 = decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_wkupidx_2 = decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_wkupidx_3 = decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_wkupidx_4 = decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_0_wkupidx_5 = decode_unit_io_macuio_3_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_valid = decode_unit_io_macuio_3_bits_srcreq_1_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_isgroup = decode_unit_io_macuio_3_bits_srcreq_1_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_iscoef = decode_unit_io_macuio_3_bits_srcreq_1_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_idx = decode_unit_io_macuio_3_bits_srcreq_1_idx; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_busy = decode_unit_io_macuio_3_bits_srcreq_1_busy; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_wkupidx_0 = decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_wkupidx_1 = decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_wkupidx_2 = decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_wkupidx_3 = decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_wkupidx_4 = decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_1_wkupidx_5 = decode_unit_io_macuio_3_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_valid = decode_unit_io_macuio_3_bits_srcreq_2_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_isgroup = decode_unit_io_macuio_3_bits_srcreq_2_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_iscoef = decode_unit_io_macuio_3_bits_srcreq_2_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_idx = decode_unit_io_macuio_3_bits_srcreq_2_idx; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_busy = decode_unit_io_macuio_3_bits_srcreq_2_busy; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_wkupidx_0 = decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_wkupidx_1 = decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_wkupidx_2 = decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_wkupidx_3 = decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_wkupidx_4 = decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_2_wkupidx_5 = decode_unit_io_macuio_3_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_valid = decode_unit_io_macuio_3_bits_srcreq_3_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_isgroup = decode_unit_io_macuio_3_bits_srcreq_3_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_iscoef = decode_unit_io_macuio_3_bits_srcreq_3_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_idx = decode_unit_io_macuio_3_bits_srcreq_3_idx; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_busy = decode_unit_io_macuio_3_bits_srcreq_3_busy; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_wkupidx_0 = decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_wkupidx_1 = decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_wkupidx_2 = decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_wkupidx_3 = decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_wkupidx_4 = decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_3_wkupidx_5 = decode_unit_io_macuio_3_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_valid = decode_unit_io_macuio_3_bits_srcreq_4_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_isgroup = decode_unit_io_macuio_3_bits_srcreq_4_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_iscoef = decode_unit_io_macuio_3_bits_srcreq_4_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_idx = decode_unit_io_macuio_3_bits_srcreq_4_idx; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_busy = decode_unit_io_macuio_3_bits_srcreq_4_busy; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_wkupidx_0 = decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_wkupidx_1 = decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_wkupidx_2 = decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_wkupidx_3 = decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_wkupidx_4 = decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_4_wkupidx_5 = decode_unit_io_macuio_3_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_valid = decode_unit_io_macuio_3_bits_srcreq_5_valid; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_isgroup = decode_unit_io_macuio_3_bits_srcreq_5_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_iscoef = decode_unit_io_macuio_3_bits_srcreq_5_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_idx = decode_unit_io_macuio_3_bits_srcreq_5_idx; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_busy = decode_unit_io_macuio_3_bits_srcreq_5_busy; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_wkupidx_0 = decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_wkupidx_1 = decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_wkupidx_2 = decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_wkupidx_3 = decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_wkupidx_4 = decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_srcreq_5_wkupidx_5 = decode_unit_io_macuio_3_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wbvld = decode_unit_io_macuio_3_bits_wbvld; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wbreq = decode_unit_io_macuio_3_bits_wbreq; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_waridx_0 = decode_unit_io_macuio_3_bits_waridx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_waridx_1 = decode_unit_io_macuio_3_bits_waridx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_waridx_2 = decode_unit_io_macuio_3_bits_waridx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_waridx_3 = decode_unit_io_macuio_3_bits_waridx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_waridx_4 = decode_unit_io_macuio_3_bits_waridx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wawidx_0 = decode_unit_io_macuio_3_bits_wawidx_0; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wawidx_1 = decode_unit_io_macuio_3_bits_wawidx_1; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wawidx_2 = decode_unit_io_macuio_3_bits_wawidx_2; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wawidx_3 = decode_unit_io_macuio_3_bits_wawidx_3; // @[dsptop.scala 171:27]
  assign mac_units_3_io_uopin_bits_wawidx_4 = decode_unit_io_macuio_3_bits_wawidx_4; // @[dsptop.scala 171:27]
  assign mac_units_3_io_rfreq_0_resp = reg_file_io_exe_rd_6_resp; // @[dsptop.scala 192:31]
  assign mac_units_3_io_rfreq_1_resp = reg_file_io_exe_rd_7_resp; // @[dsptop.scala 193:35]
  assign mac_units_3_io_raw_wkup_0_valid = mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_0_bits = mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_1_valid = mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_1_bits = mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_2_valid = mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_2_bits = mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_3_valid = mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_3_bits = mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_4_valid = mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_4_bits = mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_3_io_raw_wkup_5_valid = cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_3_io_raw_wkup_5_bits = cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_3_io_other_flop_0 = mac_units_0_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_3_io_other_flop_1 = mac_units_1_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_3_io_other_flop_2 = mac_units_2_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_3_io_other_flop_3 = mac_units_4_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_3_io_other_flop_4 = cor_unit_io_flop; // @[dsptop.scala 205:25 dsptop.scala 216:22]
  assign mac_units_3_io_coef_subch_drc_th = io_coefin_regmap_subch_drc2_coef[95:64]; // @[dsptop.scala 105:56]
  assign mac_units_3_io_coef_subch_drc_offset = {coef_subch_drc_offset_hi,coef_subch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_3_io_coef_subch_drc_drcen = io_coefin_regmap_subch_drc2_en; // @[dsptop.scala 90:25 dsptop.scala 102:24]
  assign mac_units_3_io_coef_mainch_ch0_autoloop = io_coefin_regmap_mainch_alp_en; // @[dsptop.scala 90:25 dsptop.scala 109:28]
  assign mac_units_3_io_coef_mainch_drc_th = io_coefin_regmap_mainch_drc1_coef[95:64]; // @[dsptop.scala 98:58]
  assign mac_units_3_io_coef_mainch_drc_offset = {coef_mainch_drc_offset_hi,coef_mainch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_3_io_coef_mainch_drc_drcen = io_coefin_regmap_mainch_drc1_en; // @[dsptop.scala 90:25 dsptop.scala 95:25]
  assign mac_units_4_clock = clock;
  assign mac_units_4_reset = reset;
  assign mac_units_4_io_uopin_valid = decode_unit_io_macuio_4_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_vlen = decode_unit_io_macuio_4_bits_vlen; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_select = decode_unit_io_macuio_4_bits_select; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_drc = decode_unit_io_macuio_4_bits_drc; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_pow = decode_unit_io_macuio_4_bits_pow; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_loop = decode_unit_io_macuio_4_bits_loop; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_drcgain = decode_unit_io_macuio_4_bits_drcgain; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_drcnum = decode_unit_io_macuio_4_bits_drcnum; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_valid = decode_unit_io_macuio_4_bits_srcreq_0_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_isgroup = decode_unit_io_macuio_4_bits_srcreq_0_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_iscoef = decode_unit_io_macuio_4_bits_srcreq_0_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_idx = decode_unit_io_macuio_4_bits_srcreq_0_idx; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_busy = decode_unit_io_macuio_4_bits_srcreq_0_busy; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_wkupidx_0 = decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_wkupidx_1 = decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_wkupidx_2 = decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_wkupidx_3 = decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_wkupidx_4 = decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_0_wkupidx_5 = decode_unit_io_macuio_4_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_valid = decode_unit_io_macuio_4_bits_srcreq_1_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_isgroup = decode_unit_io_macuio_4_bits_srcreq_1_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_iscoef = decode_unit_io_macuio_4_bits_srcreq_1_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_idx = decode_unit_io_macuio_4_bits_srcreq_1_idx; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_busy = decode_unit_io_macuio_4_bits_srcreq_1_busy; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_wkupidx_0 = decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_wkupidx_1 = decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_wkupidx_2 = decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_wkupidx_3 = decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_wkupidx_4 = decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_1_wkupidx_5 = decode_unit_io_macuio_4_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_valid = decode_unit_io_macuio_4_bits_srcreq_2_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_isgroup = decode_unit_io_macuio_4_bits_srcreq_2_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_iscoef = decode_unit_io_macuio_4_bits_srcreq_2_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_idx = decode_unit_io_macuio_4_bits_srcreq_2_idx; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_busy = decode_unit_io_macuio_4_bits_srcreq_2_busy; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_wkupidx_0 = decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_wkupidx_1 = decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_wkupidx_2 = decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_wkupidx_3 = decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_wkupidx_4 = decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_2_wkupidx_5 = decode_unit_io_macuio_4_bits_srcreq_2_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_valid = decode_unit_io_macuio_4_bits_srcreq_3_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_isgroup = decode_unit_io_macuio_4_bits_srcreq_3_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_iscoef = decode_unit_io_macuio_4_bits_srcreq_3_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_idx = decode_unit_io_macuio_4_bits_srcreq_3_idx; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_busy = decode_unit_io_macuio_4_bits_srcreq_3_busy; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_wkupidx_0 = decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_wkupidx_1 = decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_wkupidx_2 = decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_wkupidx_3 = decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_wkupidx_4 = decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_3_wkupidx_5 = decode_unit_io_macuio_4_bits_srcreq_3_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_valid = decode_unit_io_macuio_4_bits_srcreq_4_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_isgroup = decode_unit_io_macuio_4_bits_srcreq_4_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_iscoef = decode_unit_io_macuio_4_bits_srcreq_4_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_idx = decode_unit_io_macuio_4_bits_srcreq_4_idx; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_busy = decode_unit_io_macuio_4_bits_srcreq_4_busy; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_wkupidx_0 = decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_wkupidx_1 = decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_wkupidx_2 = decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_wkupidx_3 = decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_wkupidx_4 = decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_4_wkupidx_5 = decode_unit_io_macuio_4_bits_srcreq_4_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_valid = decode_unit_io_macuio_4_bits_srcreq_5_valid; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_isgroup = decode_unit_io_macuio_4_bits_srcreq_5_isgroup; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_iscoef = decode_unit_io_macuio_4_bits_srcreq_5_iscoef; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_idx = decode_unit_io_macuio_4_bits_srcreq_5_idx; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_busy = decode_unit_io_macuio_4_bits_srcreq_5_busy; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_wkupidx_0 = decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_wkupidx_1 = decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_wkupidx_2 = decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_wkupidx_3 = decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_wkupidx_4 = decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_srcreq_5_wkupidx_5 = decode_unit_io_macuio_4_bits_srcreq_5_wkupidx_5; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wbvld = decode_unit_io_macuio_4_bits_wbvld; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wbreq = decode_unit_io_macuio_4_bits_wbreq; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_waridx_0 = decode_unit_io_macuio_4_bits_waridx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_waridx_1 = decode_unit_io_macuio_4_bits_waridx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_waridx_2 = decode_unit_io_macuio_4_bits_waridx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_waridx_3 = decode_unit_io_macuio_4_bits_waridx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_waridx_4 = decode_unit_io_macuio_4_bits_waridx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wawidx_0 = decode_unit_io_macuio_4_bits_wawidx_0; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wawidx_1 = decode_unit_io_macuio_4_bits_wawidx_1; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wawidx_2 = decode_unit_io_macuio_4_bits_wawidx_2; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wawidx_3 = decode_unit_io_macuio_4_bits_wawidx_3; // @[dsptop.scala 171:27]
  assign mac_units_4_io_uopin_bits_wawidx_4 = decode_unit_io_macuio_4_bits_wawidx_4; // @[dsptop.scala 171:27]
  assign mac_units_4_io_rfreq_0_resp = reg_file_io_exe_rd_8_resp; // @[dsptop.scala 192:31]
  assign mac_units_4_io_rfreq_1_resp = reg_file_io_exe_rd_9_resp; // @[dsptop.scala 193:35]
  assign mac_units_4_io_raw_wkup_0_valid = mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_0_bits = mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_1_valid = mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_1_bits = mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_2_valid = mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_2_bits = mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_3_valid = mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_3_bits = mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_4_valid = mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_4_bits = mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign mac_units_4_io_raw_wkup_5_valid = cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_4_io_raw_wkup_5_bits = cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign mac_units_4_io_other_flop_0 = mac_units_0_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_4_io_other_flop_1 = mac_units_1_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_4_io_other_flop_2 = mac_units_2_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_4_io_other_flop_3 = mac_units_3_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign mac_units_4_io_other_flop_4 = cor_unit_io_flop; // @[dsptop.scala 205:25 dsptop.scala 216:22]
  assign mac_units_4_io_coef_subch_drc_th = io_coefin_regmap_subch_drc2_coef[95:64]; // @[dsptop.scala 105:56]
  assign mac_units_4_io_coef_subch_drc_offset = {coef_subch_drc_offset_hi,coef_subch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_4_io_coef_subch_drc_drcen = io_coefin_regmap_subch_drc2_en; // @[dsptop.scala 90:25 dsptop.scala 102:24]
  assign mac_units_4_io_coef_mainch_ch0_autoloop = io_coefin_regmap_mainch_alp_en; // @[dsptop.scala 90:25 dsptop.scala 109:28]
  assign mac_units_4_io_coef_mainch_drc_th = io_coefin_regmap_mainch_drc1_coef[95:64]; // @[dsptop.scala 98:58]
  assign mac_units_4_io_coef_mainch_drc_offset = {coef_mainch_drc_offset_hi,coef_mainch_drc_offset_lo}; // @[Cat.scala 30:58]
  assign mac_units_4_io_coef_mainch_drc_drcen = io_coefin_regmap_mainch_drc1_en; // @[dsptop.scala 90:25 dsptop.scala 95:25]
  assign cor_unit_clock = clock;
  assign cor_unit_reset = reset;
  assign cor_unit_io_uopin_valid = decode_unit_io_coruio_valid; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_cortype = decode_unit_io_coruio_bits_cortype; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_valid = decode_unit_io_coruio_bits_srcreq_0_valid; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_idx = decode_unit_io_coruio_bits_srcreq_0_idx; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_busy = decode_unit_io_coruio_bits_srcreq_0_busy; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_wkupidx_0 = decode_unit_io_coruio_bits_srcreq_0_wkupidx_0; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_wkupidx_1 = decode_unit_io_coruio_bits_srcreq_0_wkupidx_1; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_wkupidx_2 = decode_unit_io_coruio_bits_srcreq_0_wkupidx_2; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_wkupidx_3 = decode_unit_io_coruio_bits_srcreq_0_wkupidx_3; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_wkupidx_4 = decode_unit_io_coruio_bits_srcreq_0_wkupidx_4; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_0_wkupidx_5 = decode_unit_io_coruio_bits_srcreq_0_wkupidx_5; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_valid = decode_unit_io_coruio_bits_srcreq_1_valid; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_idx = decode_unit_io_coruio_bits_srcreq_1_idx; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_busy = decode_unit_io_coruio_bits_srcreq_1_busy; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_wkupidx_0 = decode_unit_io_coruio_bits_srcreq_1_wkupidx_0; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_wkupidx_1 = decode_unit_io_coruio_bits_srcreq_1_wkupidx_1; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_wkupidx_2 = decode_unit_io_coruio_bits_srcreq_1_wkupidx_2; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_wkupidx_3 = decode_unit_io_coruio_bits_srcreq_1_wkupidx_3; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_wkupidx_4 = decode_unit_io_coruio_bits_srcreq_1_wkupidx_4; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_srcreq_1_wkupidx_5 = decode_unit_io_coruio_bits_srcreq_1_wkupidx_5; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wbvld = decode_unit_io_coruio_bits_wbvld; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wbreq = decode_unit_io_coruio_bits_wbreq; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_waridx_0 = decode_unit_io_coruio_bits_waridx_0; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_waridx_1 = decode_unit_io_coruio_bits_waridx_1; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_waridx_2 = decode_unit_io_coruio_bits_waridx_2; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_waridx_3 = decode_unit_io_coruio_bits_waridx_3; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_waridx_4 = decode_unit_io_coruio_bits_waridx_4; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wawidx_0 = decode_unit_io_coruio_bits_wawidx_0; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wawidx_1 = decode_unit_io_coruio_bits_wawidx_1; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wawidx_2 = decode_unit_io_coruio_bits_wawidx_2; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wawidx_3 = decode_unit_io_coruio_bits_wawidx_3; // @[dsptop.scala 180:21]
  assign cor_unit_io_uopin_bits_wawidx_4 = decode_unit_io_coruio_bits_wawidx_4; // @[dsptop.scala 180:21]
  assign cor_unit_io_rfreq_0_resp = reg_file_io_exe_rd_10_resp; // @[dsptop.scala 197:36]
  assign cor_unit_io_rfreq_1_resp = reg_file_io_exe_rd_11_resp; // @[dsptop.scala 198:40]
  assign cor_unit_io_raw_wkup_0_valid = mac_units_0_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_0_bits = mac_units_0_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_1_valid = mac_units_1_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_1_bits = mac_units_1_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_2_valid = mac_units_2_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_2_bits = mac_units_2_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_3_valid = mac_units_3_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_3_bits = mac_units_3_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_4_valid = mac_units_4_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_4_bits = mac_units_4_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 209:15]
  assign cor_unit_io_raw_wkup_5_valid = cor_unit_io_fwd_wkup_valid; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign cor_unit_io_raw_wkup_5_bits = cor_unit_io_fwd_wkup_bits; // @[dsptop.scala 204:23 dsptop.scala 217:20]
  assign cor_unit_io_other_flop_0 = mac_units_0_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign cor_unit_io_other_flop_1 = mac_units_1_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign cor_unit_io_other_flop_2 = mac_units_2_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign cor_unit_io_other_flop_3 = mac_units_3_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
  assign cor_unit_io_other_flop_4 = mac_units_4_io_flop; // @[dsptop.scala 205:25 dsptop.scala 208:17]
endmodule
